library ieee;
use ieee.std_logic_1164.all;

entity eager_fork_register_block is
  port (
    clk, rst : in std_logic;
    -- inputs
    ins_valid    : in std_logic;
    outs_ready   : in std_logic;
    backpressure : in std_logic;
    -- outputs
    outs_valid : out std_logic;
    blockStop  : out std_logic
  );
end entity;

architecture arch of eager_fork_register_block is
  signal transmitValue, keepValue : std_logic;
begin
  keepValue <= (not outs_ready) and transmitValue;

  process (rst, clk)
  begin
    if (rst = '1') then
      transmitValue <= '1';
    elsif (rising_edge(clk)) then
      transmitValue <= keepValue or (not backpressure);
    end if;
  end process;

  outs_valid <= transmitValue and ins_valid;
  blockStop  <= keepValue;
end architecture;
