module mul_4_stage #(
  parameter BITWIDTH = 32
)(
  // inputs
  input  clk,
  input  ce,
  input  [BITWIDTH - 1 : 0] a,
  input  [BITWIDTH - 1 : 0] b,
  // outputs
  output [BITWIDTH - 1 : 0] p
);

  reg  [BITWIDTH - 1 : 0] a_reg;
  reg  [BITWIDTH - 1 : 0] b_reg;
  reg  [BITWIDTH - 1 : 0] q0;
  reg  [BITWIDTH - 1 : 0] q1;
  reg  [BITWIDTH - 1 : 0] q2;
  wire  [BITWIDTH - 1 : 0] mul;

  assign mul = a_reg * b_reg;

  always @(posedge clk) begin
    if (ce) begin
      a_reg <= a;
      b_reg <= b;
      q0 <= mul;
      q1 <= q0;
      q2 <= q1;
    end
  end

  assign p = q2;

endmodule


module muli #(
  parameter BITWIDTH = 32,
  parameter LATENCY = 4
)(
  // inputs
  input  clk,
  input  rst,
  input  [BITWIDTH - 1 : 0] lhs,
  input  lhs_valid,
  input  [BITWIDTH - 1 : 0] rhs,
  input  rhs_valid,
  input  result_ready,
  // outputs
  output [BITWIDTH - 1 : 0] result,
  output result_valid,
  output lhs_ready,
  output rhs_ready
);

  assert(LATENCY != 4) else $fatal("muli only supports LATENCY = 4");

  wire join_valid;
  wire oehb_ready;
  wire buff_valid;
  wire [BITWIDTH - 1 : 0] oehb_dataOut, oehb_dataIn;

  // Instantiate the join node
  join #(
    .SIZE(2)
  ) join_inputs (
    .ins_valid  ({rhs_valid, lhs_valid}),
    .outs_ready (oehb_ready             ),
    .ins_ready  ({rhs_ready, lhs_ready}  ),
    .outs_valid (join_valid             )
  );

  mul_4_stage #(
    .BITWIDTH(BITWIDTH)
  ) mul_4_stage_inst (
    .clk(clk),
    .ce(oehb_ready),
    .a(lhs),
    .b(rhs),
    .p(result)
  );

  delay_buffer #(
    .SIZE( LATENCY - 1)
  ) buff (
    .clk(clk),
    .rst(rst),
    .valid_in(join_valid),
    .ready_in(oehb_ready),
    .valid_out(buff_valid)
  );

  oehb #(
    .BITWIDTH(BITWIDTH)
  ) oehb_inst (
    .clk(clk),
    .rst(rst),
    .ins(oehb_dataIn),
    .ins_valid(buff_valid),
    .ins_ready(oehb_ready),
    .outs(oehb_dataOut),
    .outs_valid(result_valid),
    .outs_ready(result_ready)
  );


endmodule