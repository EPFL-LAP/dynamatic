library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity fork_dataless is
  generic (
    SIZE : integer
  );
  port (
    clk, rst : in std_logic;
    -- input channel
    ins_valid : in  std_logic;
    ins_ready : out std_logic;
    -- output channels
    outs_valid : out std_logic_vector(SIZE - 1 downto 0);
    outs_ready : in  std_logic_vector(SIZE - 1 downto 0)
  );
end entity;

architecture arch of fork_dataless is
  signal blockStopArray : std_logic_vector(SIZE - 1 downto 0);
  signal anyBlockStop   : std_logic;
  signal backpressure   : std_logic;
begin
  anyBlockFull : entity work.or_n generic map (SIZE)
    port map(
      blockStopArray,
      anyBlockStop
    );

  ins_ready    <= not anyBlockStop;
  backpressure <= ins_valid and anyBlockStop;

  generateBlocks : for i in SIZE - 1 downto 0 generate
    regblock : entity work.eager_fork_register_block(arch)
      port map(
        -- inputs
        clk          => clk,
        rst          => rst,
        ins_valid    => ins_valid,
        outs_ready   => outs_ready(i),
        backpressure => backpressure,
        -- outputs
        outs_valid => outs_valid(i),
        blockStop  => blockStopArray(i)
      );
  end generate;

end architecture;

entity fork_dataless_with_tag is
  generic (
    SIZE : integer
  );
  port (
    clk, rst : in std_logic;
    -- input channel
    ins_valid : in  std_logic;
    ins_spec_tag : in std_logic;
    ins_ready : out std_logic;
    -- output channels
    outs_valid : out std_logic_vector(SIZE - 1 downto 0);
    outs_spec_tag : out std_logic_vector(SIZE - 1 downto 0);
    outs_ready : in  std_logic_vector(SIZE - 1 downto 0)
  );
end entity;

architecture arch of fork_dataless_with_tag is
  signal outs : std_logic_vector(0 downto 0)
begin
  -- This is actually fork with 1-bit data
  outs_spec_tag <= outs(0);
  fork_inner : entity work.handshake_fork(arch)
    generic map(
      SIZE => SIZE,
      DATA_TYPE => 1
    )
    port map(
      clk        => clk,
      rst        => rst,
      ins => std_logic_vector(ins_spec_tag), -- todo
      ins_valid  => ins_valid,
      ins_ready  => ins_ready,
      outs => outs, -- todo
      outs_valid => outs_valid,
      outs_ready => outs_ready
    )
end architecture;
