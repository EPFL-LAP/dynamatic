library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity kernel_3mm is
  port (
    A_loadData : in std_logic_vector(31 downto 0);
    B_loadData : in std_logic_vector(31 downto 0);
    C_loadData : in std_logic_vector(31 downto 0);
    D_loadData : in std_logic_vector(31 downto 0);
    E_loadData : in std_logic_vector(31 downto 0);
    F_loadData : in std_logic_vector(31 downto 0);
    G_loadData : in std_logic_vector(31 downto 0);
    A_start_valid : in std_logic;
    B_start_valid : in std_logic;
    C_start_valid : in std_logic;
    D_start_valid : in std_logic;
    E_start_valid : in std_logic;
    F_start_valid : in std_logic;
    G_start_valid : in std_logic;
    start_valid : in std_logic;
    clk : in std_logic;
    rst : in std_logic;
    A_end_ready : in std_logic;
    B_end_ready : in std_logic;
    C_end_ready : in std_logic;
    D_end_ready : in std_logic;
    E_end_ready : in std_logic;
    F_end_ready : in std_logic;
    G_end_ready : in std_logic;
    end_ready : in std_logic;
    A_start_ready : out std_logic;
    B_start_ready : out std_logic;
    C_start_ready : out std_logic;
    D_start_ready : out std_logic;
    E_start_ready : out std_logic;
    F_start_ready : out std_logic;
    G_start_ready : out std_logic;
    start_ready : out std_logic;
    A_end_valid : out std_logic;
    B_end_valid : out std_logic;
    C_end_valid : out std_logic;
    D_end_valid : out std_logic;
    E_end_valid : out std_logic;
    F_end_valid : out std_logic;
    G_end_valid : out std_logic;
    end_valid : out std_logic;
    A_loadEn : out std_logic;
    A_loadAddr : out std_logic_vector(6 downto 0);
    A_storeEn : out std_logic;
    A_storeAddr : out std_logic_vector(6 downto 0);
    A_storeData : out std_logic_vector(31 downto 0);
    B_loadEn : out std_logic;
    B_loadAddr : out std_logic_vector(6 downto 0);
    B_storeEn : out std_logic;
    B_storeAddr : out std_logic_vector(6 downto 0);
    B_storeData : out std_logic_vector(31 downto 0);
    C_loadEn : out std_logic;
    C_loadAddr : out std_logic_vector(6 downto 0);
    C_storeEn : out std_logic;
    C_storeAddr : out std_logic_vector(6 downto 0);
    C_storeData : out std_logic_vector(31 downto 0);
    D_loadEn : out std_logic;
    D_loadAddr : out std_logic_vector(6 downto 0);
    D_storeEn : out std_logic;
    D_storeAddr : out std_logic_vector(6 downto 0);
    D_storeData : out std_logic_vector(31 downto 0);
    E_loadEn : out std_logic;
    E_loadAddr : out std_logic_vector(6 downto 0);
    E_storeEn : out std_logic;
    E_storeAddr : out std_logic_vector(6 downto 0);
    E_storeData : out std_logic_vector(31 downto 0);
    F_loadEn : out std_logic;
    F_loadAddr : out std_logic_vector(6 downto 0);
    F_storeEn : out std_logic;
    F_storeAddr : out std_logic_vector(6 downto 0);
    F_storeData : out std_logic_vector(31 downto 0);
    G_loadEn : out std_logic;
    G_loadAddr : out std_logic_vector(6 downto 0);
    G_storeEn : out std_logic;
    G_storeAddr : out std_logic_vector(6 downto 0);
    G_storeData : out std_logic_vector(31 downto 0)
  );
end entity;

architecture behavioral of kernel_3mm is

  signal fork0_outs_0_valid : std_logic;
  signal fork0_outs_0_ready : std_logic;
  signal fork0_outs_1_valid : std_logic;
  signal fork0_outs_1_ready : std_logic;
  signal fork0_outs_2_valid : std_logic;
  signal fork0_outs_2_ready : std_logic;
  signal fork0_outs_3_valid : std_logic;
  signal fork0_outs_3_ready : std_logic;
  signal fork0_outs_4_valid : std_logic;
  signal fork0_outs_4_ready : std_logic;
  signal fork0_outs_5_valid : std_logic;
  signal fork0_outs_5_ready : std_logic;
  signal mem_controller4_stDone_0_valid : std_logic;
  signal mem_controller4_stDone_0_ready : std_logic;
  signal mem_controller4_ldData_0 : std_logic_vector(31 downto 0);
  signal mem_controller4_ldData_0_valid : std_logic;
  signal mem_controller4_ldData_0_ready : std_logic;
  signal mem_controller4_stDone_1_valid : std_logic;
  signal mem_controller4_stDone_1_ready : std_logic;
  signal mem_controller4_memEnd_valid : std_logic;
  signal mem_controller4_memEnd_ready : std_logic;
  signal mem_controller4_loadEn : std_logic;
  signal mem_controller4_loadAddr : std_logic_vector(6 downto 0);
  signal mem_controller4_storeEn : std_logic;
  signal mem_controller4_storeAddr : std_logic_vector(6 downto 0);
  signal mem_controller4_storeData : std_logic_vector(31 downto 0);
  signal mem_controller5_stDone_0_valid : std_logic;
  signal mem_controller5_stDone_0_ready : std_logic;
  signal mem_controller5_ldData_0 : std_logic_vector(31 downto 0);
  signal mem_controller5_ldData_0_valid : std_logic;
  signal mem_controller5_ldData_0_ready : std_logic;
  signal mem_controller5_stDone_1_valid : std_logic;
  signal mem_controller5_stDone_1_ready : std_logic;
  signal mem_controller5_ldData_1 : std_logic_vector(31 downto 0);
  signal mem_controller5_ldData_1_valid : std_logic;
  signal mem_controller5_ldData_1_ready : std_logic;
  signal mem_controller5_memEnd_valid : std_logic;
  signal mem_controller5_memEnd_ready : std_logic;
  signal mem_controller5_loadEn : std_logic;
  signal mem_controller5_loadAddr : std_logic_vector(6 downto 0);
  signal mem_controller5_storeEn : std_logic;
  signal mem_controller5_storeAddr : std_logic_vector(6 downto 0);
  signal mem_controller5_storeData : std_logic_vector(31 downto 0);
  signal mem_controller6_stDone_0_valid : std_logic;
  signal mem_controller6_stDone_0_ready : std_logic;
  signal mem_controller6_ldData_0 : std_logic_vector(31 downto 0);
  signal mem_controller6_ldData_0_valid : std_logic;
  signal mem_controller6_ldData_0_ready : std_logic;
  signal mem_controller6_stDone_1_valid : std_logic;
  signal mem_controller6_stDone_1_ready : std_logic;
  signal mem_controller6_ldData_1 : std_logic_vector(31 downto 0);
  signal mem_controller6_ldData_1_valid : std_logic;
  signal mem_controller6_ldData_1_ready : std_logic;
  signal mem_controller6_memEnd_valid : std_logic;
  signal mem_controller6_memEnd_ready : std_logic;
  signal mem_controller6_loadEn : std_logic;
  signal mem_controller6_loadAddr : std_logic_vector(6 downto 0);
  signal mem_controller6_storeEn : std_logic;
  signal mem_controller6_storeAddr : std_logic_vector(6 downto 0);
  signal mem_controller6_storeData : std_logic_vector(31 downto 0);
  signal mem_controller7_ldData_0 : std_logic_vector(31 downto 0);
  signal mem_controller7_ldData_0_valid : std_logic;
  signal mem_controller7_ldData_0_ready : std_logic;
  signal mem_controller7_memEnd_valid : std_logic;
  signal mem_controller7_memEnd_ready : std_logic;
  signal mem_controller7_loadEn : std_logic;
  signal mem_controller7_loadAddr : std_logic_vector(6 downto 0);
  signal mem_controller7_storeEn : std_logic;
  signal mem_controller7_storeAddr : std_logic_vector(6 downto 0);
  signal mem_controller7_storeData : std_logic_vector(31 downto 0);
  signal mem_controller8_ldData_0 : std_logic_vector(31 downto 0);
  signal mem_controller8_ldData_0_valid : std_logic;
  signal mem_controller8_ldData_0_ready : std_logic;
  signal mem_controller8_memEnd_valid : std_logic;
  signal mem_controller8_memEnd_ready : std_logic;
  signal mem_controller8_loadEn : std_logic;
  signal mem_controller8_loadAddr : std_logic_vector(6 downto 0);
  signal mem_controller8_storeEn : std_logic;
  signal mem_controller8_storeAddr : std_logic_vector(6 downto 0);
  signal mem_controller8_storeData : std_logic_vector(31 downto 0);
  signal mem_controller9_ldData_0 : std_logic_vector(31 downto 0);
  signal mem_controller9_ldData_0_valid : std_logic;
  signal mem_controller9_ldData_0_ready : std_logic;
  signal mem_controller9_memEnd_valid : std_logic;
  signal mem_controller9_memEnd_ready : std_logic;
  signal mem_controller9_loadEn : std_logic;
  signal mem_controller9_loadAddr : std_logic_vector(6 downto 0);
  signal mem_controller9_storeEn : std_logic;
  signal mem_controller9_storeAddr : std_logic_vector(6 downto 0);
  signal mem_controller9_storeData : std_logic_vector(31 downto 0);
  signal mem_controller10_ldData_0 : std_logic_vector(31 downto 0);
  signal mem_controller10_ldData_0_valid : std_logic;
  signal mem_controller10_ldData_0_ready : std_logic;
  signal mem_controller10_memEnd_valid : std_logic;
  signal mem_controller10_memEnd_ready : std_logic;
  signal mem_controller10_loadEn : std_logic;
  signal mem_controller10_loadAddr : std_logic_vector(6 downto 0);
  signal mem_controller10_storeEn : std_logic;
  signal mem_controller10_storeAddr : std_logic_vector(6 downto 0);
  signal mem_controller10_storeData : std_logic_vector(31 downto 0);
  signal constant45_outs : std_logic_vector(0 downto 0);
  signal constant45_outs_valid : std_logic;
  signal constant45_outs_ready : std_logic;
  signal extsi53_outs : std_logic_vector(4 downto 0);
  signal extsi53_outs_valid : std_logic;
  signal extsi53_outs_ready : std_logic;
  signal mux22_outs_valid : std_logic;
  signal mux22_outs_ready : std_logic;
  signal init0_outs : std_logic_vector(0 downto 0);
  signal init0_outs_valid : std_logic;
  signal init0_outs_ready : std_logic;
  signal mux0_outs : std_logic_vector(4 downto 0);
  signal mux0_outs_valid : std_logic;
  signal mux0_outs_ready : std_logic;
  signal control_merge0_outs_valid : std_logic;
  signal control_merge0_outs_ready : std_logic;
  signal control_merge0_index : std_logic_vector(0 downto 0);
  signal control_merge0_index_valid : std_logic;
  signal control_merge0_index_ready : std_logic;
  signal fork1_outs_0_valid : std_logic;
  signal fork1_outs_0_ready : std_logic;
  signal fork1_outs_1_valid : std_logic;
  signal fork1_outs_1_ready : std_logic;
  signal constant46_outs : std_logic_vector(0 downto 0);
  signal constant46_outs_valid : std_logic;
  signal constant46_outs_ready : std_logic;
  signal extsi52_outs : std_logic_vector(4 downto 0);
  signal extsi52_outs_valid : std_logic;
  signal extsi52_outs_ready : std_logic;
  signal buffer8_outs : std_logic_vector(4 downto 0);
  signal buffer8_outs_valid : std_logic;
  signal buffer8_outs_ready : std_logic;
  signal buffer6_outs_valid : std_logic;
  signal buffer6_outs_ready : std_logic;
  signal mux27_outs_valid : std_logic;
  signal mux27_outs_ready : std_logic;
  signal init5_outs : std_logic_vector(0 downto 0);
  signal init5_outs_valid : std_logic;
  signal init5_outs_ready : std_logic;
  signal buffer7_outs : std_logic_vector(0 downto 0);
  signal buffer7_outs_valid : std_logic;
  signal buffer7_outs_ready : std_logic;
  signal mux1_outs : std_logic_vector(4 downto 0);
  signal mux1_outs_valid : std_logic;
  signal mux1_outs_ready : std_logic;
  signal buffer11_outs : std_logic_vector(4 downto 0);
  signal buffer11_outs_valid : std_logic;
  signal buffer11_outs_ready : std_logic;
  signal fork2_outs_0 : std_logic_vector(4 downto 0);
  signal fork2_outs_0_valid : std_logic;
  signal fork2_outs_0_ready : std_logic;
  signal fork2_outs_1 : std_logic_vector(4 downto 0);
  signal fork2_outs_1_valid : std_logic;
  signal fork2_outs_1_ready : std_logic;
  signal extsi54_outs : std_logic_vector(6 downto 0);
  signal extsi54_outs_valid : std_logic;
  signal extsi54_outs_ready : std_logic;
  signal mux2_outs : std_logic_vector(4 downto 0);
  signal mux2_outs_valid : std_logic;
  signal mux2_outs_ready : std_logic;
  signal buffer12_outs : std_logic_vector(4 downto 0);
  signal buffer12_outs_valid : std_logic;
  signal buffer12_outs_ready : std_logic;
  signal buffer13_outs : std_logic_vector(4 downto 0);
  signal buffer13_outs_valid : std_logic;
  signal buffer13_outs_ready : std_logic;
  signal fork3_outs_0 : std_logic_vector(4 downto 0);
  signal fork3_outs_0_valid : std_logic;
  signal fork3_outs_0_ready : std_logic;
  signal fork3_outs_1 : std_logic_vector(4 downto 0);
  signal fork3_outs_1_valid : std_logic;
  signal fork3_outs_1_ready : std_logic;
  signal extsi55_outs : std_logic_vector(31 downto 0);
  signal extsi55_outs_valid : std_logic;
  signal extsi55_outs_ready : std_logic;
  signal fork4_outs_0 : std_logic_vector(31 downto 0);
  signal fork4_outs_0_valid : std_logic;
  signal fork4_outs_0_ready : std_logic;
  signal fork4_outs_1 : std_logic_vector(31 downto 0);
  signal fork4_outs_1_valid : std_logic;
  signal fork4_outs_1_ready : std_logic;
  signal control_merge1_outs_valid : std_logic;
  signal control_merge1_outs_ready : std_logic;
  signal control_merge1_index : std_logic_vector(0 downto 0);
  signal control_merge1_index_valid : std_logic;
  signal control_merge1_index_ready : std_logic;
  signal fork5_outs_0 : std_logic_vector(0 downto 0);
  signal fork5_outs_0_valid : std_logic;
  signal fork5_outs_0_ready : std_logic;
  signal fork5_outs_1 : std_logic_vector(0 downto 0);
  signal fork5_outs_1_valid : std_logic;
  signal fork5_outs_1_ready : std_logic;
  signal fork6_outs_0_valid : std_logic;
  signal fork6_outs_0_ready : std_logic;
  signal fork6_outs_1_valid : std_logic;
  signal fork6_outs_1_ready : std_logic;
  signal fork6_outs_2_valid : std_logic;
  signal fork6_outs_2_ready : std_logic;
  signal constant47_outs : std_logic_vector(1 downto 0);
  signal constant47_outs_valid : std_logic;
  signal constant47_outs_ready : std_logic;
  signal extsi2_outs : std_logic_vector(31 downto 0);
  signal extsi2_outs_valid : std_logic;
  signal extsi2_outs_ready : std_logic;
  signal constant48_outs : std_logic_vector(0 downto 0);
  signal constant48_outs_valid : std_logic;
  signal constant48_outs_ready : std_logic;
  signal fork7_outs_0 : std_logic_vector(0 downto 0);
  signal fork7_outs_0_valid : std_logic;
  signal fork7_outs_0_ready : std_logic;
  signal fork7_outs_1 : std_logic_vector(0 downto 0);
  signal fork7_outs_1_valid : std_logic;
  signal fork7_outs_1_ready : std_logic;
  signal extsi4_outs : std_logic_vector(31 downto 0);
  signal extsi4_outs_valid : std_logic;
  signal extsi4_outs_ready : std_logic;
  signal source0_outs_valid : std_logic;
  signal source0_outs_ready : std_logic;
  signal constant49_outs : std_logic_vector(1 downto 0);
  signal constant49_outs_valid : std_logic;
  signal constant49_outs_ready : std_logic;
  signal extsi5_outs : std_logic_vector(31 downto 0);
  signal extsi5_outs_valid : std_logic;
  signal extsi5_outs_ready : std_logic;
  signal source1_outs_valid : std_logic;
  signal source1_outs_ready : std_logic;
  signal constant50_outs : std_logic_vector(2 downto 0);
  signal constant50_outs_valid : std_logic;
  signal constant50_outs_ready : std_logic;
  signal extsi6_outs : std_logic_vector(31 downto 0);
  signal extsi6_outs_valid : std_logic;
  signal extsi6_outs_ready : std_logic;
  signal shli0_result : std_logic_vector(31 downto 0);
  signal shli0_result_valid : std_logic;
  signal shli0_result_ready : std_logic;
  signal buffer14_outs : std_logic_vector(31 downto 0);
  signal buffer14_outs_valid : std_logic;
  signal buffer14_outs_ready : std_logic;
  signal trunci0_outs : std_logic_vector(6 downto 0);
  signal trunci0_outs_valid : std_logic;
  signal trunci0_outs_ready : std_logic;
  signal shli1_result : std_logic_vector(31 downto 0);
  signal shli1_result_valid : std_logic;
  signal shli1_result_ready : std_logic;
  signal buffer15_outs : std_logic_vector(31 downto 0);
  signal buffer15_outs_valid : std_logic;
  signal buffer15_outs_ready : std_logic;
  signal trunci1_outs : std_logic_vector(6 downto 0);
  signal trunci1_outs_valid : std_logic;
  signal trunci1_outs_ready : std_logic;
  signal addi27_result : std_logic_vector(6 downto 0);
  signal addi27_result_valid : std_logic;
  signal addi27_result_ready : std_logic;
  signal buffer16_outs : std_logic_vector(6 downto 0);
  signal buffer16_outs_valid : std_logic;
  signal buffer16_outs_ready : std_logic;
  signal addi3_result : std_logic_vector(6 downto 0);
  signal addi3_result_valid : std_logic;
  signal addi3_result_ready : std_logic;
  signal buffer0_outs_valid : std_logic;
  signal buffer0_outs_ready : std_logic;
  signal fork8_outs_0_valid : std_logic;
  signal fork8_outs_0_ready : std_logic;
  signal fork8_outs_1_valid : std_logic;
  signal fork8_outs_1_ready : std_logic;
  signal buffer17_outs : std_logic_vector(6 downto 0);
  signal buffer17_outs_valid : std_logic;
  signal buffer17_outs_ready : std_logic;
  signal store0_addrOut : std_logic_vector(6 downto 0);
  signal store0_addrOut_valid : std_logic;
  signal store0_addrOut_ready : std_logic;
  signal store0_dataToMem : std_logic_vector(31 downto 0);
  signal store0_dataToMem_valid : std_logic;
  signal store0_dataToMem_ready : std_logic;
  signal store0_doneOut_valid : std_logic;
  signal store0_doneOut_ready : std_logic;
  signal extsi51_outs : std_logic_vector(4 downto 0);
  signal extsi51_outs_valid : std_logic;
  signal extsi51_outs_ready : std_logic;
  signal buffer65_outs_valid : std_logic;
  signal buffer65_outs_ready : std_logic;
  signal cond_br116_trueOut_valid : std_logic;
  signal cond_br116_trueOut_ready : std_logic;
  signal cond_br116_falseOut_valid : std_logic;
  signal cond_br116_falseOut_ready : std_logic;
  signal buffer18_outs : std_logic_vector(0 downto 0);
  signal buffer18_outs_valid : std_logic;
  signal buffer18_outs_ready : std_logic;
  signal cond_br117_trueOut_valid : std_logic;
  signal cond_br117_trueOut_ready : std_logic;
  signal cond_br117_falseOut_valid : std_logic;
  signal cond_br117_falseOut_ready : std_logic;
  signal buffer19_outs : std_logic_vector(0 downto 0);
  signal buffer19_outs_valid : std_logic;
  signal buffer19_outs_ready : std_logic;
  signal init10_outs : std_logic_vector(0 downto 0);
  signal init10_outs_valid : std_logic;
  signal init10_outs_ready : std_logic;
  signal fork9_outs_0 : std_logic_vector(0 downto 0);
  signal fork9_outs_0_valid : std_logic;
  signal fork9_outs_0_ready : std_logic;
  signal fork9_outs_1 : std_logic_vector(0 downto 0);
  signal fork9_outs_1_valid : std_logic;
  signal fork9_outs_1_ready : std_logic;
  signal mux28_outs_valid : std_logic;
  signal mux28_outs_ready : std_logic;
  signal buffer21_outs : std_logic_vector(0 downto 0);
  signal buffer21_outs_valid : std_logic;
  signal buffer21_outs_ready : std_logic;
  signal buffer20_outs_valid : std_logic;
  signal buffer20_outs_ready : std_logic;
  signal buffer23_outs_valid : std_logic;
  signal buffer23_outs_ready : std_logic;
  signal fork10_outs_0_valid : std_logic;
  signal fork10_outs_0_ready : std_logic;
  signal fork10_outs_1_valid : std_logic;
  signal fork10_outs_1_ready : std_logic;
  signal fork10_outs_2_valid : std_logic;
  signal fork10_outs_2_ready : std_logic;
  signal buffer9_outs_valid : std_logic;
  signal buffer9_outs_ready : std_logic;
  signal buffer10_outs_valid : std_logic;
  signal buffer10_outs_ready : std_logic;
  signal mux31_outs_valid : std_logic;
  signal mux31_outs_ready : std_logic;
  signal buffer22_outs : std_logic_vector(0 downto 0);
  signal buffer22_outs_valid : std_logic;
  signal buffer22_outs_ready : std_logic;
  signal mux3_outs : std_logic_vector(4 downto 0);
  signal mux3_outs_valid : std_logic;
  signal mux3_outs_ready : std_logic;
  signal buffer26_outs : std_logic_vector(4 downto 0);
  signal buffer26_outs_valid : std_logic;
  signal buffer26_outs_ready : std_logic;
  signal buffer27_outs : std_logic_vector(4 downto 0);
  signal buffer27_outs_valid : std_logic;
  signal buffer27_outs_ready : std_logic;
  signal fork11_outs_0 : std_logic_vector(4 downto 0);
  signal fork11_outs_0_valid : std_logic;
  signal fork11_outs_0_ready : std_logic;
  signal fork11_outs_1 : std_logic_vector(4 downto 0);
  signal fork11_outs_1_valid : std_logic;
  signal fork11_outs_1_ready : std_logic;
  signal fork11_outs_2 : std_logic_vector(4 downto 0);
  signal fork11_outs_2_valid : std_logic;
  signal fork11_outs_2_ready : std_logic;
  signal extsi56_outs : std_logic_vector(6 downto 0);
  signal extsi56_outs_valid : std_logic;
  signal extsi56_outs_ready : std_logic;
  signal buffer24_outs : std_logic_vector(4 downto 0);
  signal buffer24_outs_valid : std_logic;
  signal buffer24_outs_ready : std_logic;
  signal extsi57_outs : std_logic_vector(5 downto 0);
  signal extsi57_outs_valid : std_logic;
  signal extsi57_outs_ready : std_logic;
  signal extsi58_outs : std_logic_vector(31 downto 0);
  signal extsi58_outs_valid : std_logic;
  signal extsi58_outs_ready : std_logic;
  signal fork12_outs_0 : std_logic_vector(31 downto 0);
  signal fork12_outs_0_valid : std_logic;
  signal fork12_outs_0_ready : std_logic;
  signal fork12_outs_1 : std_logic_vector(31 downto 0);
  signal fork12_outs_1_valid : std_logic;
  signal fork12_outs_1_ready : std_logic;
  signal mux4_outs : std_logic_vector(4 downto 0);
  signal mux4_outs_valid : std_logic;
  signal mux4_outs_ready : std_logic;
  signal buffer28_outs : std_logic_vector(4 downto 0);
  signal buffer28_outs_valid : std_logic;
  signal buffer28_outs_ready : std_logic;
  signal buffer29_outs : std_logic_vector(4 downto 0);
  signal buffer29_outs_valid : std_logic;
  signal buffer29_outs_ready : std_logic;
  signal fork13_outs_0 : std_logic_vector(4 downto 0);
  signal fork13_outs_0_valid : std_logic;
  signal fork13_outs_0_ready : std_logic;
  signal fork13_outs_1 : std_logic_vector(4 downto 0);
  signal fork13_outs_1_valid : std_logic;
  signal fork13_outs_1_ready : std_logic;
  signal extsi59_outs : std_logic_vector(31 downto 0);
  signal extsi59_outs_valid : std_logic;
  signal extsi59_outs_ready : std_logic;
  signal fork14_outs_0 : std_logic_vector(31 downto 0);
  signal fork14_outs_0_valid : std_logic;
  signal fork14_outs_0_ready : std_logic;
  signal fork14_outs_1 : std_logic_vector(31 downto 0);
  signal fork14_outs_1_valid : std_logic;
  signal fork14_outs_1_ready : std_logic;
  signal fork14_outs_2 : std_logic_vector(31 downto 0);
  signal fork14_outs_2_valid : std_logic;
  signal fork14_outs_2_ready : std_logic;
  signal fork14_outs_3 : std_logic_vector(31 downto 0);
  signal fork14_outs_3_valid : std_logic;
  signal fork14_outs_3_ready : std_logic;
  signal fork14_outs_4 : std_logic_vector(31 downto 0);
  signal fork14_outs_4_valid : std_logic;
  signal fork14_outs_4_ready : std_logic;
  signal fork14_outs_5 : std_logic_vector(31 downto 0);
  signal fork14_outs_5_valid : std_logic;
  signal fork14_outs_5_ready : std_logic;
  signal mux5_outs : std_logic_vector(4 downto 0);
  signal mux5_outs_valid : std_logic;
  signal mux5_outs_ready : std_logic;
  signal buffer31_outs : std_logic_vector(4 downto 0);
  signal buffer31_outs_valid : std_logic;
  signal buffer31_outs_ready : std_logic;
  signal buffer34_outs : std_logic_vector(4 downto 0);
  signal buffer34_outs_valid : std_logic;
  signal buffer34_outs_ready : std_logic;
  signal fork15_outs_0 : std_logic_vector(4 downto 0);
  signal fork15_outs_0_valid : std_logic;
  signal fork15_outs_0_ready : std_logic;
  signal fork15_outs_1 : std_logic_vector(4 downto 0);
  signal fork15_outs_1_valid : std_logic;
  signal fork15_outs_1_ready : std_logic;
  signal fork15_outs_2 : std_logic_vector(4 downto 0);
  signal fork15_outs_2_valid : std_logic;
  signal fork15_outs_2_ready : std_logic;
  signal extsi60_outs : std_logic_vector(6 downto 0);
  signal extsi60_outs_valid : std_logic;
  signal extsi60_outs_ready : std_logic;
  signal buffer30_outs : std_logic_vector(4 downto 0);
  signal buffer30_outs_valid : std_logic;
  signal buffer30_outs_ready : std_logic;
  signal extsi61_outs : std_logic_vector(31 downto 0);
  signal extsi61_outs_valid : std_logic;
  signal extsi61_outs_ready : std_logic;
  signal fork16_outs_0 : std_logic_vector(31 downto 0);
  signal fork16_outs_0_valid : std_logic;
  signal fork16_outs_0_ready : std_logic;
  signal fork16_outs_1 : std_logic_vector(31 downto 0);
  signal fork16_outs_1_valid : std_logic;
  signal fork16_outs_1_ready : std_logic;
  signal control_merge2_outs_valid : std_logic;
  signal control_merge2_outs_ready : std_logic;
  signal control_merge2_index : std_logic_vector(0 downto 0);
  signal control_merge2_index_valid : std_logic;
  signal control_merge2_index_ready : std_logic;
  signal fork17_outs_0 : std_logic_vector(0 downto 0);
  signal fork17_outs_0_valid : std_logic;
  signal fork17_outs_0_ready : std_logic;
  signal fork17_outs_1 : std_logic_vector(0 downto 0);
  signal fork17_outs_1_valid : std_logic;
  signal fork17_outs_1_ready : std_logic;
  signal fork17_outs_2 : std_logic_vector(0 downto 0);
  signal fork17_outs_2_valid : std_logic;
  signal fork17_outs_2_ready : std_logic;
  signal fork18_outs_0_valid : std_logic;
  signal fork18_outs_0_ready : std_logic;
  signal fork18_outs_1_valid : std_logic;
  signal fork18_outs_1_ready : std_logic;
  signal constant51_outs : std_logic_vector(1 downto 0);
  signal constant51_outs_valid : std_logic;
  signal constant51_outs_ready : std_logic;
  signal extsi7_outs : std_logic_vector(31 downto 0);
  signal extsi7_outs_valid : std_logic;
  signal extsi7_outs_ready : std_logic;
  signal source2_outs_valid : std_logic;
  signal source2_outs_ready : std_logic;
  signal constant52_outs : std_logic_vector(4 downto 0);
  signal constant52_outs_valid : std_logic;
  signal constant52_outs_ready : std_logic;
  signal extsi62_outs : std_logic_vector(5 downto 0);
  signal extsi62_outs_valid : std_logic;
  signal extsi62_outs_ready : std_logic;
  signal source3_outs_valid : std_logic;
  signal source3_outs_ready : std_logic;
  signal constant53_outs : std_logic_vector(1 downto 0);
  signal constant53_outs_valid : std_logic;
  signal constant53_outs_ready : std_logic;
  signal fork19_outs_0 : std_logic_vector(1 downto 0);
  signal fork19_outs_0_valid : std_logic;
  signal fork19_outs_0_ready : std_logic;
  signal fork19_outs_1 : std_logic_vector(1 downto 0);
  signal fork19_outs_1_valid : std_logic;
  signal fork19_outs_1_ready : std_logic;
  signal extsi63_outs : std_logic_vector(5 downto 0);
  signal extsi63_outs_valid : std_logic;
  signal extsi63_outs_ready : std_logic;
  signal buffer32_outs : std_logic_vector(1 downto 0);
  signal buffer32_outs_valid : std_logic;
  signal buffer32_outs_ready : std_logic;
  signal extsi9_outs : std_logic_vector(31 downto 0);
  signal extsi9_outs_valid : std_logic;
  signal extsi9_outs_ready : std_logic;
  signal buffer33_outs : std_logic_vector(1 downto 0);
  signal buffer33_outs_valid : std_logic;
  signal buffer33_outs_ready : std_logic;
  signal fork20_outs_0 : std_logic_vector(31 downto 0);
  signal fork20_outs_0_valid : std_logic;
  signal fork20_outs_0_ready : std_logic;
  signal fork20_outs_1 : std_logic_vector(31 downto 0);
  signal fork20_outs_1_valid : std_logic;
  signal fork20_outs_1_ready : std_logic;
  signal fork20_outs_2 : std_logic_vector(31 downto 0);
  signal fork20_outs_2_valid : std_logic;
  signal fork20_outs_2_ready : std_logic;
  signal fork20_outs_3 : std_logic_vector(31 downto 0);
  signal fork20_outs_3_valid : std_logic;
  signal fork20_outs_3_ready : std_logic;
  signal source4_outs_valid : std_logic;
  signal source4_outs_ready : std_logic;
  signal constant54_outs : std_logic_vector(2 downto 0);
  signal constant54_outs_valid : std_logic;
  signal constant54_outs_ready : std_logic;
  signal extsi10_outs : std_logic_vector(31 downto 0);
  signal extsi10_outs_valid : std_logic;
  signal extsi10_outs_ready : std_logic;
  signal fork21_outs_0 : std_logic_vector(31 downto 0);
  signal fork21_outs_0_valid : std_logic;
  signal fork21_outs_0_ready : std_logic;
  signal fork21_outs_1 : std_logic_vector(31 downto 0);
  signal fork21_outs_1_valid : std_logic;
  signal fork21_outs_1_ready : std_logic;
  signal fork21_outs_2 : std_logic_vector(31 downto 0);
  signal fork21_outs_2_valid : std_logic;
  signal fork21_outs_2_ready : std_logic;
  signal fork21_outs_3 : std_logic_vector(31 downto 0);
  signal fork21_outs_3_valid : std_logic;
  signal fork21_outs_3_ready : std_logic;
  signal shli2_result : std_logic_vector(31 downto 0);
  signal shli2_result_valid : std_logic;
  signal shli2_result_ready : std_logic;
  signal buffer35_outs : std_logic_vector(31 downto 0);
  signal buffer35_outs_valid : std_logic;
  signal buffer35_outs_ready : std_logic;
  signal buffer38_outs : std_logic_vector(31 downto 0);
  signal buffer38_outs_valid : std_logic;
  signal buffer38_outs_ready : std_logic;
  signal trunci2_outs : std_logic_vector(6 downto 0);
  signal trunci2_outs_valid : std_logic;
  signal trunci2_outs_ready : std_logic;
  signal shli3_result : std_logic_vector(31 downto 0);
  signal shli3_result_valid : std_logic;
  signal shli3_result_ready : std_logic;
  signal buffer37_outs : std_logic_vector(31 downto 0);
  signal buffer37_outs_valid : std_logic;
  signal buffer37_outs_ready : std_logic;
  signal buffer40_outs : std_logic_vector(31 downto 0);
  signal buffer40_outs_valid : std_logic;
  signal buffer40_outs_ready : std_logic;
  signal trunci3_outs : std_logic_vector(6 downto 0);
  signal trunci3_outs_valid : std_logic;
  signal trunci3_outs_ready : std_logic;
  signal addi28_result : std_logic_vector(6 downto 0);
  signal addi28_result_valid : std_logic;
  signal addi28_result_ready : std_logic;
  signal buffer52_outs : std_logic_vector(6 downto 0);
  signal buffer52_outs_valid : std_logic;
  signal buffer52_outs_ready : std_logic;
  signal addi4_result : std_logic_vector(6 downto 0);
  signal addi4_result_valid : std_logic;
  signal addi4_result_ready : std_logic;
  signal load0_addrOut : std_logic_vector(6 downto 0);
  signal load0_addrOut_valid : std_logic;
  signal load0_addrOut_ready : std_logic;
  signal load0_dataOut : std_logic_vector(31 downto 0);
  signal load0_dataOut_valid : std_logic;
  signal load0_dataOut_ready : std_logic;
  signal shli4_result : std_logic_vector(31 downto 0);
  signal shli4_result_valid : std_logic;
  signal shli4_result_ready : std_logic;
  signal buffer39_outs : std_logic_vector(31 downto 0);
  signal buffer39_outs_valid : std_logic;
  signal buffer39_outs_ready : std_logic;
  signal buffer53_outs : std_logic_vector(31 downto 0);
  signal buffer53_outs_valid : std_logic;
  signal buffer53_outs_ready : std_logic;
  signal trunci4_outs : std_logic_vector(6 downto 0);
  signal trunci4_outs_valid : std_logic;
  signal trunci4_outs_ready : std_logic;
  signal shli5_result : std_logic_vector(31 downto 0);
  signal shli5_result_valid : std_logic;
  signal shli5_result_ready : std_logic;
  signal buffer41_outs : std_logic_vector(31 downto 0);
  signal buffer41_outs_valid : std_logic;
  signal buffer41_outs_ready : std_logic;
  signal buffer54_outs : std_logic_vector(31 downto 0);
  signal buffer54_outs_valid : std_logic;
  signal buffer54_outs_ready : std_logic;
  signal trunci5_outs : std_logic_vector(6 downto 0);
  signal trunci5_outs_valid : std_logic;
  signal trunci5_outs_ready : std_logic;
  signal addi29_result : std_logic_vector(6 downto 0);
  signal addi29_result_valid : std_logic;
  signal addi29_result_ready : std_logic;
  signal buffer56_outs : std_logic_vector(6 downto 0);
  signal buffer56_outs_valid : std_logic;
  signal buffer56_outs_ready : std_logic;
  signal addi5_result : std_logic_vector(6 downto 0);
  signal addi5_result_valid : std_logic;
  signal addi5_result_ready : std_logic;
  signal load1_addrOut : std_logic_vector(6 downto 0);
  signal load1_addrOut_valid : std_logic;
  signal load1_addrOut_ready : std_logic;
  signal load1_dataOut : std_logic_vector(31 downto 0);
  signal load1_dataOut_valid : std_logic;
  signal load1_dataOut_ready : std_logic;
  signal muli0_result : std_logic_vector(31 downto 0);
  signal muli0_result_valid : std_logic;
  signal muli0_result_ready : std_logic;
  signal shli6_result : std_logic_vector(31 downto 0);
  signal shli6_result_valid : std_logic;
  signal shli6_result_ready : std_logic;
  signal buffer42_outs : std_logic_vector(31 downto 0);
  signal buffer42_outs_valid : std_logic;
  signal buffer42_outs_ready : std_logic;
  signal buffer43_outs : std_logic_vector(31 downto 0);
  signal buffer43_outs_valid : std_logic;
  signal buffer43_outs_ready : std_logic;
  signal shli7_result : std_logic_vector(31 downto 0);
  signal shli7_result_valid : std_logic;
  signal shli7_result_ready : std_logic;
  signal buffer44_outs : std_logic_vector(31 downto 0);
  signal buffer44_outs_valid : std_logic;
  signal buffer44_outs_ready : std_logic;
  signal buffer45_outs : std_logic_vector(31 downto 0);
  signal buffer45_outs_valid : std_logic;
  signal buffer45_outs_ready : std_logic;
  signal buffer57_outs : std_logic_vector(31 downto 0);
  signal buffer57_outs_valid : std_logic;
  signal buffer57_outs_ready : std_logic;
  signal buffer58_outs : std_logic_vector(31 downto 0);
  signal buffer58_outs_valid : std_logic;
  signal buffer58_outs_ready : std_logic;
  signal addi30_result : std_logic_vector(31 downto 0);
  signal addi30_result_valid : std_logic;
  signal addi30_result_ready : std_logic;
  signal buffer61_outs : std_logic_vector(31 downto 0);
  signal buffer61_outs_valid : std_logic;
  signal buffer61_outs_ready : std_logic;
  signal addi6_result : std_logic_vector(31 downto 0);
  signal addi6_result_valid : std_logic;
  signal addi6_result_ready : std_logic;
  signal buffer46_outs : std_logic_vector(31 downto 0);
  signal buffer46_outs_valid : std_logic;
  signal buffer46_outs_ready : std_logic;
  signal buffer25_outs_valid : std_logic;
  signal buffer25_outs_ready : std_logic;
  signal gate0_outs : std_logic_vector(31 downto 0);
  signal gate0_outs_valid : std_logic;
  signal gate0_outs_ready : std_logic;
  signal trunci6_outs : std_logic_vector(6 downto 0);
  signal trunci6_outs_valid : std_logic;
  signal trunci6_outs_ready : std_logic;
  signal load2_addrOut : std_logic_vector(6 downto 0);
  signal load2_addrOut_valid : std_logic;
  signal load2_addrOut_ready : std_logic;
  signal load2_dataOut : std_logic_vector(31 downto 0);
  signal load2_dataOut_valid : std_logic;
  signal load2_dataOut_ready : std_logic;
  signal addi0_result : std_logic_vector(31 downto 0);
  signal addi0_result_valid : std_logic;
  signal addi0_result_ready : std_logic;
  signal shli8_result : std_logic_vector(31 downto 0);
  signal shli8_result_valid : std_logic;
  signal shli8_result_ready : std_logic;
  signal buffer47_outs : std_logic_vector(31 downto 0);
  signal buffer47_outs_valid : std_logic;
  signal buffer47_outs_ready : std_logic;
  signal buffer48_outs : std_logic_vector(31 downto 0);
  signal buffer48_outs_valid : std_logic;
  signal buffer48_outs_ready : std_logic;
  signal shli9_result : std_logic_vector(31 downto 0);
  signal shli9_result_valid : std_logic;
  signal shli9_result_ready : std_logic;
  signal buffer49_outs : std_logic_vector(31 downto 0);
  signal buffer49_outs_valid : std_logic;
  signal buffer49_outs_ready : std_logic;
  signal buffer50_outs : std_logic_vector(31 downto 0);
  signal buffer50_outs_valid : std_logic;
  signal buffer50_outs_ready : std_logic;
  signal buffer62_outs : std_logic_vector(31 downto 0);
  signal buffer62_outs_valid : std_logic;
  signal buffer62_outs_ready : std_logic;
  signal buffer63_outs : std_logic_vector(31 downto 0);
  signal buffer63_outs_valid : std_logic;
  signal buffer63_outs_ready : std_logic;
  signal addi31_result : std_logic_vector(31 downto 0);
  signal addi31_result_valid : std_logic;
  signal addi31_result_ready : std_logic;
  signal buffer64_outs : std_logic_vector(31 downto 0);
  signal buffer64_outs_valid : std_logic;
  signal buffer64_outs_ready : std_logic;
  signal addi7_result : std_logic_vector(31 downto 0);
  signal addi7_result_valid : std_logic;
  signal addi7_result_ready : std_logic;
  signal buffer51_outs : std_logic_vector(31 downto 0);
  signal buffer51_outs_valid : std_logic;
  signal buffer51_outs_ready : std_logic;
  signal buffer1_outs_valid : std_logic;
  signal buffer1_outs_ready : std_logic;
  signal gate1_outs : std_logic_vector(31 downto 0);
  signal gate1_outs_valid : std_logic;
  signal gate1_outs_ready : std_logic;
  signal trunci7_outs : std_logic_vector(6 downto 0);
  signal trunci7_outs_valid : std_logic;
  signal trunci7_outs_ready : std_logic;
  signal store1_addrOut : std_logic_vector(6 downto 0);
  signal store1_addrOut_valid : std_logic;
  signal store1_addrOut_ready : std_logic;
  signal store1_dataToMem : std_logic_vector(31 downto 0);
  signal store1_dataToMem_valid : std_logic;
  signal store1_dataToMem_ready : std_logic;
  signal store1_doneOut_valid : std_logic;
  signal store1_doneOut_ready : std_logic;
  signal addi18_result : std_logic_vector(5 downto 0);
  signal addi18_result_valid : std_logic;
  signal addi18_result_ready : std_logic;
  signal buffer67_outs : std_logic_vector(5 downto 0);
  signal buffer67_outs_valid : std_logic;
  signal buffer67_outs_ready : std_logic;
  signal fork22_outs_0 : std_logic_vector(5 downto 0);
  signal fork22_outs_0_valid : std_logic;
  signal fork22_outs_0_ready : std_logic;
  signal fork22_outs_1 : std_logic_vector(5 downto 0);
  signal fork22_outs_1_valid : std_logic;
  signal fork22_outs_1_ready : std_logic;
  signal trunci8_outs : std_logic_vector(4 downto 0);
  signal trunci8_outs_valid : std_logic;
  signal trunci8_outs_ready : std_logic;
  signal cmpi0_result : std_logic_vector(0 downto 0);
  signal cmpi0_result_valid : std_logic;
  signal cmpi0_result_ready : std_logic;
  signal buffer68_outs : std_logic_vector(0 downto 0);
  signal buffer68_outs_valid : std_logic;
  signal buffer68_outs_ready : std_logic;
  signal fork23_outs_0 : std_logic_vector(0 downto 0);
  signal fork23_outs_0_valid : std_logic;
  signal fork23_outs_0_ready : std_logic;
  signal fork23_outs_1 : std_logic_vector(0 downto 0);
  signal fork23_outs_1_valid : std_logic;
  signal fork23_outs_1_ready : std_logic;
  signal fork23_outs_2 : std_logic_vector(0 downto 0);
  signal fork23_outs_2_valid : std_logic;
  signal fork23_outs_2_ready : std_logic;
  signal fork23_outs_3 : std_logic_vector(0 downto 0);
  signal fork23_outs_3_valid : std_logic;
  signal fork23_outs_3_ready : std_logic;
  signal fork23_outs_4 : std_logic_vector(0 downto 0);
  signal fork23_outs_4_valid : std_logic;
  signal fork23_outs_4_ready : std_logic;
  signal fork23_outs_5 : std_logic_vector(0 downto 0);
  signal fork23_outs_5_valid : std_logic;
  signal fork23_outs_5_ready : std_logic;
  signal fork23_outs_6 : std_logic_vector(0 downto 0);
  signal fork23_outs_6_valid : std_logic;
  signal fork23_outs_6_ready : std_logic;
  signal cond_br9_trueOut : std_logic_vector(4 downto 0);
  signal cond_br9_trueOut_valid : std_logic;
  signal cond_br9_trueOut_ready : std_logic;
  signal cond_br9_falseOut : std_logic_vector(4 downto 0);
  signal cond_br9_falseOut_valid : std_logic;
  signal cond_br9_falseOut_ready : std_logic;
  signal cond_br10_trueOut : std_logic_vector(4 downto 0);
  signal cond_br10_trueOut_valid : std_logic;
  signal cond_br10_trueOut_ready : std_logic;
  signal cond_br10_falseOut : std_logic_vector(4 downto 0);
  signal cond_br10_falseOut_valid : std_logic;
  signal cond_br10_falseOut_ready : std_logic;
  signal buffer55_outs : std_logic_vector(0 downto 0);
  signal buffer55_outs_valid : std_logic;
  signal buffer55_outs_ready : std_logic;
  signal cond_br11_trueOut : std_logic_vector(4 downto 0);
  signal cond_br11_trueOut_valid : std_logic;
  signal cond_br11_trueOut_ready : std_logic;
  signal cond_br11_falseOut : std_logic_vector(4 downto 0);
  signal cond_br11_falseOut_valid : std_logic;
  signal cond_br11_falseOut_ready : std_logic;
  signal buffer36_outs_valid : std_logic;
  signal buffer36_outs_ready : std_logic;
  signal cond_br12_trueOut_valid : std_logic;
  signal cond_br12_trueOut_ready : std_logic;
  signal cond_br12_falseOut_valid : std_logic;
  signal cond_br12_falseOut_ready : std_logic;
  signal buffer59_outs : std_logic_vector(0 downto 0);
  signal buffer59_outs_valid : std_logic;
  signal buffer59_outs_ready : std_logic;
  signal cond_br118_trueOut_valid : std_logic;
  signal cond_br118_trueOut_ready : std_logic;
  signal cond_br118_falseOut_valid : std_logic;
  signal cond_br118_falseOut_ready : std_logic;
  signal buffer60_outs : std_logic_vector(0 downto 0);
  signal buffer60_outs_valid : std_logic;
  signal buffer60_outs_ready : std_logic;
  signal cond_br119_trueOut_valid : std_logic;
  signal cond_br119_trueOut_ready : std_logic;
  signal cond_br119_falseOut_valid : std_logic;
  signal cond_br119_falseOut_ready : std_logic;
  signal extsi64_outs : std_logic_vector(5 downto 0);
  signal extsi64_outs_valid : std_logic;
  signal extsi64_outs_ready : std_logic;
  signal source5_outs_valid : std_logic;
  signal source5_outs_ready : std_logic;
  signal constant55_outs : std_logic_vector(4 downto 0);
  signal constant55_outs_valid : std_logic;
  signal constant55_outs_ready : std_logic;
  signal extsi65_outs : std_logic_vector(5 downto 0);
  signal extsi65_outs_valid : std_logic;
  signal extsi65_outs_ready : std_logic;
  signal source6_outs_valid : std_logic;
  signal source6_outs_ready : std_logic;
  signal constant56_outs : std_logic_vector(1 downto 0);
  signal constant56_outs_valid : std_logic;
  signal constant56_outs_ready : std_logic;
  signal extsi66_outs : std_logic_vector(5 downto 0);
  signal extsi66_outs_valid : std_logic;
  signal extsi66_outs_ready : std_logic;
  signal addi19_result : std_logic_vector(5 downto 0);
  signal addi19_result_valid : std_logic;
  signal addi19_result_ready : std_logic;
  signal buffer69_outs : std_logic_vector(5 downto 0);
  signal buffer69_outs_valid : std_logic;
  signal buffer69_outs_ready : std_logic;
  signal fork24_outs_0 : std_logic_vector(5 downto 0);
  signal fork24_outs_0_valid : std_logic;
  signal fork24_outs_0_ready : std_logic;
  signal fork24_outs_1 : std_logic_vector(5 downto 0);
  signal fork24_outs_1_valid : std_logic;
  signal fork24_outs_1_ready : std_logic;
  signal trunci9_outs : std_logic_vector(4 downto 0);
  signal trunci9_outs_valid : std_logic;
  signal trunci9_outs_ready : std_logic;
  signal cmpi1_result : std_logic_vector(0 downto 0);
  signal cmpi1_result_valid : std_logic;
  signal cmpi1_result_ready : std_logic;
  signal buffer70_outs : std_logic_vector(0 downto 0);
  signal buffer70_outs_valid : std_logic;
  signal buffer70_outs_ready : std_logic;
  signal fork25_outs_0 : std_logic_vector(0 downto 0);
  signal fork25_outs_0_valid : std_logic;
  signal fork25_outs_0_ready : std_logic;
  signal fork25_outs_1 : std_logic_vector(0 downto 0);
  signal fork25_outs_1_valid : std_logic;
  signal fork25_outs_1_ready : std_logic;
  signal fork25_outs_2 : std_logic_vector(0 downto 0);
  signal fork25_outs_2_valid : std_logic;
  signal fork25_outs_2_ready : std_logic;
  signal fork25_outs_3 : std_logic_vector(0 downto 0);
  signal fork25_outs_3_valid : std_logic;
  signal fork25_outs_3_ready : std_logic;
  signal fork25_outs_4 : std_logic_vector(0 downto 0);
  signal fork25_outs_4_valid : std_logic;
  signal fork25_outs_4_ready : std_logic;
  signal fork25_outs_5 : std_logic_vector(0 downto 0);
  signal fork25_outs_5_valid : std_logic;
  signal fork25_outs_5_ready : std_logic;
  signal cond_br13_trueOut : std_logic_vector(4 downto 0);
  signal cond_br13_trueOut_valid : std_logic;
  signal cond_br13_trueOut_ready : std_logic;
  signal cond_br13_falseOut : std_logic_vector(4 downto 0);
  signal cond_br13_falseOut_valid : std_logic;
  signal cond_br13_falseOut_ready : std_logic;
  signal cond_br14_trueOut : std_logic_vector(4 downto 0);
  signal cond_br14_trueOut_valid : std_logic;
  signal cond_br14_trueOut_ready : std_logic;
  signal cond_br14_falseOut : std_logic_vector(4 downto 0);
  signal cond_br14_falseOut_valid : std_logic;
  signal cond_br14_falseOut_ready : std_logic;
  signal cond_br15_trueOut_valid : std_logic;
  signal cond_br15_trueOut_ready : std_logic;
  signal cond_br15_falseOut_valid : std_logic;
  signal cond_br15_falseOut_ready : std_logic;
  signal buffer66_outs : std_logic_vector(0 downto 0);
  signal buffer66_outs_valid : std_logic;
  signal buffer66_outs_ready : std_logic;
  signal cond_br120_trueOut_valid : std_logic;
  signal cond_br120_trueOut_ready : std_logic;
  signal cond_br120_falseOut_valid : std_logic;
  signal cond_br120_falseOut_ready : std_logic;
  signal cond_br121_trueOut_valid : std_logic;
  signal cond_br121_trueOut_ready : std_logic;
  signal cond_br121_falseOut_valid : std_logic;
  signal cond_br121_falseOut_ready : std_logic;
  signal buffer71_outs : std_logic_vector(4 downto 0);
  signal buffer71_outs_valid : std_logic;
  signal buffer71_outs_ready : std_logic;
  signal extsi67_outs : std_logic_vector(5 downto 0);
  signal extsi67_outs_valid : std_logic;
  signal extsi67_outs_ready : std_logic;
  signal fork26_outs_0_valid : std_logic;
  signal fork26_outs_0_ready : std_logic;
  signal fork26_outs_1_valid : std_logic;
  signal fork26_outs_1_ready : std_logic;
  signal constant57_outs : std_logic_vector(0 downto 0);
  signal constant57_outs_valid : std_logic;
  signal constant57_outs_ready : std_logic;
  signal source7_outs_valid : std_logic;
  signal source7_outs_ready : std_logic;
  signal constant58_outs : std_logic_vector(4 downto 0);
  signal constant58_outs_valid : std_logic;
  signal constant58_outs_ready : std_logic;
  signal extsi68_outs : std_logic_vector(5 downto 0);
  signal extsi68_outs_valid : std_logic;
  signal extsi68_outs_ready : std_logic;
  signal source8_outs_valid : std_logic;
  signal source8_outs_ready : std_logic;
  signal constant59_outs : std_logic_vector(1 downto 0);
  signal constant59_outs_valid : std_logic;
  signal constant59_outs_ready : std_logic;
  signal extsi69_outs : std_logic_vector(5 downto 0);
  signal extsi69_outs_valid : std_logic;
  signal extsi69_outs_ready : std_logic;
  signal addi20_result : std_logic_vector(5 downto 0);
  signal addi20_result_valid : std_logic;
  signal addi20_result_ready : std_logic;
  signal buffer72_outs : std_logic_vector(5 downto 0);
  signal buffer72_outs_valid : std_logic;
  signal buffer72_outs_ready : std_logic;
  signal fork27_outs_0 : std_logic_vector(5 downto 0);
  signal fork27_outs_0_valid : std_logic;
  signal fork27_outs_0_ready : std_logic;
  signal fork27_outs_1 : std_logic_vector(5 downto 0);
  signal fork27_outs_1_valid : std_logic;
  signal fork27_outs_1_ready : std_logic;
  signal trunci10_outs : std_logic_vector(4 downto 0);
  signal trunci10_outs_valid : std_logic;
  signal trunci10_outs_ready : std_logic;
  signal cmpi2_result : std_logic_vector(0 downto 0);
  signal cmpi2_result_valid : std_logic;
  signal cmpi2_result_ready : std_logic;
  signal buffer73_outs : std_logic_vector(0 downto 0);
  signal buffer73_outs_valid : std_logic;
  signal buffer73_outs_ready : std_logic;
  signal fork28_outs_0 : std_logic_vector(0 downto 0);
  signal fork28_outs_0_valid : std_logic;
  signal fork28_outs_0_ready : std_logic;
  signal fork28_outs_1 : std_logic_vector(0 downto 0);
  signal fork28_outs_1_valid : std_logic;
  signal fork28_outs_1_ready : std_logic;
  signal fork28_outs_2 : std_logic_vector(0 downto 0);
  signal fork28_outs_2_valid : std_logic;
  signal fork28_outs_2_ready : std_logic;
  signal fork28_outs_3 : std_logic_vector(0 downto 0);
  signal fork28_outs_3_valid : std_logic;
  signal fork28_outs_3_ready : std_logic;
  signal fork28_outs_4 : std_logic_vector(0 downto 0);
  signal fork28_outs_4_valid : std_logic;
  signal fork28_outs_4_ready : std_logic;
  signal fork28_outs_5 : std_logic_vector(0 downto 0);
  signal fork28_outs_5_valid : std_logic;
  signal fork28_outs_5_ready : std_logic;
  signal cond_br16_trueOut : std_logic_vector(4 downto 0);
  signal cond_br16_trueOut_valid : std_logic;
  signal cond_br16_trueOut_ready : std_logic;
  signal cond_br16_falseOut : std_logic_vector(4 downto 0);
  signal cond_br16_falseOut_valid : std_logic;
  signal cond_br16_falseOut_ready : std_logic;
  signal cond_br17_trueOut_valid : std_logic;
  signal cond_br17_trueOut_ready : std_logic;
  signal cond_br17_falseOut_valid : std_logic;
  signal cond_br17_falseOut_ready : std_logic;
  signal cond_br18_trueOut : std_logic_vector(0 downto 0);
  signal cond_br18_trueOut_valid : std_logic;
  signal cond_br18_trueOut_ready : std_logic;
  signal cond_br18_falseOut : std_logic_vector(0 downto 0);
  signal cond_br18_falseOut_valid : std_logic;
  signal cond_br18_falseOut_ready : std_logic;
  signal extsi50_outs : std_logic_vector(4 downto 0);
  signal extsi50_outs_valid : std_logic;
  signal extsi50_outs_ready : std_logic;
  signal mux35_outs_valid : std_logic;
  signal mux35_outs_ready : std_logic;
  signal init14_outs : std_logic_vector(0 downto 0);
  signal init14_outs_valid : std_logic;
  signal init14_outs_ready : std_logic;
  signal mux6_outs : std_logic_vector(4 downto 0);
  signal mux6_outs_valid : std_logic;
  signal mux6_outs_ready : std_logic;
  signal control_merge5_outs_valid : std_logic;
  signal control_merge5_outs_ready : std_logic;
  signal control_merge5_index : std_logic_vector(0 downto 0);
  signal control_merge5_index_valid : std_logic;
  signal control_merge5_index_ready : std_logic;
  signal fork29_outs_0_valid : std_logic;
  signal fork29_outs_0_ready : std_logic;
  signal fork29_outs_1_valid : std_logic;
  signal fork29_outs_1_ready : std_logic;
  signal constant60_outs : std_logic_vector(0 downto 0);
  signal constant60_outs_valid : std_logic;
  signal constant60_outs_ready : std_logic;
  signal extsi49_outs : std_logic_vector(4 downto 0);
  signal extsi49_outs_valid : std_logic;
  signal extsi49_outs_ready : std_logic;
  signal buffer75_outs : std_logic_vector(4 downto 0);
  signal buffer75_outs_valid : std_logic;
  signal buffer75_outs_ready : std_logic;
  signal buffer74_outs_valid : std_logic;
  signal buffer74_outs_ready : std_logic;
  signal mux40_outs_valid : std_logic;
  signal mux40_outs_ready : std_logic;
  signal init19_outs : std_logic_vector(0 downto 0);
  signal init19_outs_valid : std_logic;
  signal init19_outs_ready : std_logic;
  signal mux7_outs : std_logic_vector(4 downto 0);
  signal mux7_outs_valid : std_logic;
  signal mux7_outs_ready : std_logic;
  signal buffer78_outs : std_logic_vector(4 downto 0);
  signal buffer78_outs_valid : std_logic;
  signal buffer78_outs_ready : std_logic;
  signal fork30_outs_0 : std_logic_vector(4 downto 0);
  signal fork30_outs_0_valid : std_logic;
  signal fork30_outs_0_ready : std_logic;
  signal fork30_outs_1 : std_logic_vector(4 downto 0);
  signal fork30_outs_1_valid : std_logic;
  signal fork30_outs_1_ready : std_logic;
  signal extsi70_outs : std_logic_vector(6 downto 0);
  signal extsi70_outs_valid : std_logic;
  signal extsi70_outs_ready : std_logic;
  signal mux8_outs : std_logic_vector(4 downto 0);
  signal mux8_outs_valid : std_logic;
  signal mux8_outs_ready : std_logic;
  signal buffer79_outs : std_logic_vector(4 downto 0);
  signal buffer79_outs_valid : std_logic;
  signal buffer79_outs_ready : std_logic;
  signal buffer80_outs : std_logic_vector(4 downto 0);
  signal buffer80_outs_valid : std_logic;
  signal buffer80_outs_ready : std_logic;
  signal fork31_outs_0 : std_logic_vector(4 downto 0);
  signal fork31_outs_0_valid : std_logic;
  signal fork31_outs_0_ready : std_logic;
  signal fork31_outs_1 : std_logic_vector(4 downto 0);
  signal fork31_outs_1_valid : std_logic;
  signal fork31_outs_1_ready : std_logic;
  signal extsi71_outs : std_logic_vector(31 downto 0);
  signal extsi71_outs_valid : std_logic;
  signal extsi71_outs_ready : std_logic;
  signal fork32_outs_0 : std_logic_vector(31 downto 0);
  signal fork32_outs_0_valid : std_logic;
  signal fork32_outs_0_ready : std_logic;
  signal fork32_outs_1 : std_logic_vector(31 downto 0);
  signal fork32_outs_1_valid : std_logic;
  signal fork32_outs_1_ready : std_logic;
  signal control_merge6_outs_valid : std_logic;
  signal control_merge6_outs_ready : std_logic;
  signal control_merge6_index : std_logic_vector(0 downto 0);
  signal control_merge6_index_valid : std_logic;
  signal control_merge6_index_ready : std_logic;
  signal fork33_outs_0 : std_logic_vector(0 downto 0);
  signal fork33_outs_0_valid : std_logic;
  signal fork33_outs_0_ready : std_logic;
  signal fork33_outs_1 : std_logic_vector(0 downto 0);
  signal fork33_outs_1_valid : std_logic;
  signal fork33_outs_1_ready : std_logic;
  signal fork34_outs_0_valid : std_logic;
  signal fork34_outs_0_ready : std_logic;
  signal fork34_outs_1_valid : std_logic;
  signal fork34_outs_1_ready : std_logic;
  signal fork34_outs_2_valid : std_logic;
  signal fork34_outs_2_ready : std_logic;
  signal constant61_outs : std_logic_vector(1 downto 0);
  signal constant61_outs_valid : std_logic;
  signal constant61_outs_ready : std_logic;
  signal extsi17_outs : std_logic_vector(31 downto 0);
  signal extsi17_outs_valid : std_logic;
  signal extsi17_outs_ready : std_logic;
  signal constant62_outs : std_logic_vector(0 downto 0);
  signal constant62_outs_valid : std_logic;
  signal constant62_outs_ready : std_logic;
  signal fork35_outs_0 : std_logic_vector(0 downto 0);
  signal fork35_outs_0_valid : std_logic;
  signal fork35_outs_0_ready : std_logic;
  signal fork35_outs_1 : std_logic_vector(0 downto 0);
  signal fork35_outs_1_valid : std_logic;
  signal fork35_outs_1_ready : std_logic;
  signal extsi19_outs : std_logic_vector(31 downto 0);
  signal extsi19_outs_valid : std_logic;
  signal extsi19_outs_ready : std_logic;
  signal source9_outs_valid : std_logic;
  signal source9_outs_ready : std_logic;
  signal constant63_outs : std_logic_vector(1 downto 0);
  signal constant63_outs_valid : std_logic;
  signal constant63_outs_ready : std_logic;
  signal extsi20_outs : std_logic_vector(31 downto 0);
  signal extsi20_outs_valid : std_logic;
  signal extsi20_outs_ready : std_logic;
  signal source10_outs_valid : std_logic;
  signal source10_outs_ready : std_logic;
  signal constant64_outs : std_logic_vector(2 downto 0);
  signal constant64_outs_valid : std_logic;
  signal constant64_outs_ready : std_logic;
  signal extsi21_outs : std_logic_vector(31 downto 0);
  signal extsi21_outs_valid : std_logic;
  signal extsi21_outs_ready : std_logic;
  signal shli10_result : std_logic_vector(31 downto 0);
  signal shli10_result_valid : std_logic;
  signal shli10_result_ready : std_logic;
  signal buffer81_outs : std_logic_vector(31 downto 0);
  signal buffer81_outs_valid : std_logic;
  signal buffer81_outs_ready : std_logic;
  signal trunci11_outs : std_logic_vector(6 downto 0);
  signal trunci11_outs_valid : std_logic;
  signal trunci11_outs_ready : std_logic;
  signal shli11_result : std_logic_vector(31 downto 0);
  signal shli11_result_valid : std_logic;
  signal shli11_result_ready : std_logic;
  signal buffer82_outs : std_logic_vector(31 downto 0);
  signal buffer82_outs_valid : std_logic;
  signal buffer82_outs_ready : std_logic;
  signal trunci12_outs : std_logic_vector(6 downto 0);
  signal trunci12_outs_valid : std_logic;
  signal trunci12_outs_ready : std_logic;
  signal addi32_result : std_logic_vector(6 downto 0);
  signal addi32_result_valid : std_logic;
  signal addi32_result_ready : std_logic;
  signal buffer83_outs : std_logic_vector(6 downto 0);
  signal buffer83_outs_valid : std_logic;
  signal buffer83_outs_ready : std_logic;
  signal addi8_result : std_logic_vector(6 downto 0);
  signal addi8_result_valid : std_logic;
  signal addi8_result_ready : std_logic;
  signal buffer2_outs_valid : std_logic;
  signal buffer2_outs_ready : std_logic;
  signal fork36_outs_0_valid : std_logic;
  signal fork36_outs_0_ready : std_logic;
  signal fork36_outs_1_valid : std_logic;
  signal fork36_outs_1_ready : std_logic;
  signal buffer84_outs : std_logic_vector(6 downto 0);
  signal buffer84_outs_valid : std_logic;
  signal buffer84_outs_ready : std_logic;
  signal store2_addrOut : std_logic_vector(6 downto 0);
  signal store2_addrOut_valid : std_logic;
  signal store2_addrOut_ready : std_logic;
  signal store2_dataToMem : std_logic_vector(31 downto 0);
  signal store2_dataToMem_valid : std_logic;
  signal store2_dataToMem_ready : std_logic;
  signal store2_doneOut_valid : std_logic;
  signal store2_doneOut_ready : std_logic;
  signal extsi48_outs : std_logic_vector(4 downto 0);
  signal extsi48_outs_valid : std_logic;
  signal extsi48_outs_ready : std_logic;
  signal cond_br122_trueOut_valid : std_logic;
  signal cond_br122_trueOut_ready : std_logic;
  signal cond_br122_falseOut_valid : std_logic;
  signal cond_br122_falseOut_ready : std_logic;
  signal buffer86_outs : std_logic_vector(0 downto 0);
  signal buffer86_outs_valid : std_logic;
  signal buffer86_outs_ready : std_logic;
  signal buffer126_outs_valid : std_logic;
  signal buffer126_outs_ready : std_logic;
  signal cond_br123_trueOut_valid : std_logic;
  signal cond_br123_trueOut_ready : std_logic;
  signal cond_br123_falseOut_valid : std_logic;
  signal cond_br123_falseOut_ready : std_logic;
  signal buffer87_outs : std_logic_vector(0 downto 0);
  signal buffer87_outs_valid : std_logic;
  signal buffer87_outs_ready : std_logic;
  signal init24_outs : std_logic_vector(0 downto 0);
  signal init24_outs_valid : std_logic;
  signal init24_outs_ready : std_logic;
  signal fork37_outs_0 : std_logic_vector(0 downto 0);
  signal fork37_outs_0_valid : std_logic;
  signal fork37_outs_0_ready : std_logic;
  signal fork37_outs_1 : std_logic_vector(0 downto 0);
  signal fork37_outs_1_valid : std_logic;
  signal fork37_outs_1_ready : std_logic;
  signal mux42_outs_valid : std_logic;
  signal mux42_outs_ready : std_logic;
  signal buffer89_outs : std_logic_vector(0 downto 0);
  signal buffer89_outs_valid : std_logic;
  signal buffer89_outs_ready : std_logic;
  signal buffer85_outs_valid : std_logic;
  signal buffer85_outs_ready : std_logic;
  signal buffer88_outs_valid : std_logic;
  signal buffer88_outs_ready : std_logic;
  signal fork38_outs_0_valid : std_logic;
  signal fork38_outs_0_ready : std_logic;
  signal fork38_outs_1_valid : std_logic;
  signal fork38_outs_1_ready : std_logic;
  signal fork38_outs_2_valid : std_logic;
  signal fork38_outs_2_ready : std_logic;
  signal buffer76_outs_valid : std_logic;
  signal buffer76_outs_ready : std_logic;
  signal buffer77_outs_valid : std_logic;
  signal buffer77_outs_ready : std_logic;
  signal mux45_outs_valid : std_logic;
  signal mux45_outs_ready : std_logic;
  signal buffer90_outs : std_logic_vector(0 downto 0);
  signal buffer90_outs_valid : std_logic;
  signal buffer90_outs_ready : std_logic;
  signal mux9_outs : std_logic_vector(4 downto 0);
  signal mux9_outs_valid : std_logic;
  signal mux9_outs_ready : std_logic;
  signal buffer92_outs : std_logic_vector(4 downto 0);
  signal buffer92_outs_valid : std_logic;
  signal buffer92_outs_ready : std_logic;
  signal buffer93_outs : std_logic_vector(4 downto 0);
  signal buffer93_outs_valid : std_logic;
  signal buffer93_outs_ready : std_logic;
  signal fork39_outs_0 : std_logic_vector(4 downto 0);
  signal fork39_outs_0_valid : std_logic;
  signal fork39_outs_0_ready : std_logic;
  signal fork39_outs_1 : std_logic_vector(4 downto 0);
  signal fork39_outs_1_valid : std_logic;
  signal fork39_outs_1_ready : std_logic;
  signal fork39_outs_2 : std_logic_vector(4 downto 0);
  signal fork39_outs_2_valid : std_logic;
  signal fork39_outs_2_ready : std_logic;
  signal extsi72_outs : std_logic_vector(6 downto 0);
  signal extsi72_outs_valid : std_logic;
  signal extsi72_outs_ready : std_logic;
  signal extsi73_outs : std_logic_vector(5 downto 0);
  signal extsi73_outs_valid : std_logic;
  signal extsi73_outs_ready : std_logic;
  signal extsi74_outs : std_logic_vector(31 downto 0);
  signal extsi74_outs_valid : std_logic;
  signal extsi74_outs_ready : std_logic;
  signal fork40_outs_0 : std_logic_vector(31 downto 0);
  signal fork40_outs_0_valid : std_logic;
  signal fork40_outs_0_ready : std_logic;
  signal fork40_outs_1 : std_logic_vector(31 downto 0);
  signal fork40_outs_1_valid : std_logic;
  signal fork40_outs_1_ready : std_logic;
  signal mux10_outs : std_logic_vector(4 downto 0);
  signal mux10_outs_valid : std_logic;
  signal mux10_outs_ready : std_logic;
  signal buffer94_outs : std_logic_vector(4 downto 0);
  signal buffer94_outs_valid : std_logic;
  signal buffer94_outs_ready : std_logic;
  signal buffer95_outs : std_logic_vector(4 downto 0);
  signal buffer95_outs_valid : std_logic;
  signal buffer95_outs_ready : std_logic;
  signal fork41_outs_0 : std_logic_vector(4 downto 0);
  signal fork41_outs_0_valid : std_logic;
  signal fork41_outs_0_ready : std_logic;
  signal fork41_outs_1 : std_logic_vector(4 downto 0);
  signal fork41_outs_1_valid : std_logic;
  signal fork41_outs_1_ready : std_logic;
  signal extsi75_outs : std_logic_vector(31 downto 0);
  signal extsi75_outs_valid : std_logic;
  signal extsi75_outs_ready : std_logic;
  signal fork42_outs_0 : std_logic_vector(31 downto 0);
  signal fork42_outs_0_valid : std_logic;
  signal fork42_outs_0_ready : std_logic;
  signal fork42_outs_1 : std_logic_vector(31 downto 0);
  signal fork42_outs_1_valid : std_logic;
  signal fork42_outs_1_ready : std_logic;
  signal fork42_outs_2 : std_logic_vector(31 downto 0);
  signal fork42_outs_2_valid : std_logic;
  signal fork42_outs_2_ready : std_logic;
  signal fork42_outs_3 : std_logic_vector(31 downto 0);
  signal fork42_outs_3_valid : std_logic;
  signal fork42_outs_3_ready : std_logic;
  signal fork42_outs_4 : std_logic_vector(31 downto 0);
  signal fork42_outs_4_valid : std_logic;
  signal fork42_outs_4_ready : std_logic;
  signal fork42_outs_5 : std_logic_vector(31 downto 0);
  signal fork42_outs_5_valid : std_logic;
  signal fork42_outs_5_ready : std_logic;
  signal mux11_outs : std_logic_vector(4 downto 0);
  signal mux11_outs_valid : std_logic;
  signal mux11_outs_ready : std_logic;
  signal buffer97_outs : std_logic_vector(0 downto 0);
  signal buffer97_outs_valid : std_logic;
  signal buffer97_outs_ready : std_logic;
  signal buffer96_outs : std_logic_vector(4 downto 0);
  signal buffer96_outs_valid : std_logic;
  signal buffer96_outs_ready : std_logic;
  signal buffer98_outs : std_logic_vector(4 downto 0);
  signal buffer98_outs_valid : std_logic;
  signal buffer98_outs_ready : std_logic;
  signal fork43_outs_0 : std_logic_vector(4 downto 0);
  signal fork43_outs_0_valid : std_logic;
  signal fork43_outs_0_ready : std_logic;
  signal fork43_outs_1 : std_logic_vector(4 downto 0);
  signal fork43_outs_1_valid : std_logic;
  signal fork43_outs_1_ready : std_logic;
  signal fork43_outs_2 : std_logic_vector(4 downto 0);
  signal fork43_outs_2_valid : std_logic;
  signal fork43_outs_2_ready : std_logic;
  signal extsi76_outs : std_logic_vector(6 downto 0);
  signal extsi76_outs_valid : std_logic;
  signal extsi76_outs_ready : std_logic;
  signal extsi77_outs : std_logic_vector(31 downto 0);
  signal extsi77_outs_valid : std_logic;
  signal extsi77_outs_ready : std_logic;
  signal buffer99_outs : std_logic_vector(4 downto 0);
  signal buffer99_outs_valid : std_logic;
  signal buffer99_outs_ready : std_logic;
  signal fork44_outs_0 : std_logic_vector(31 downto 0);
  signal fork44_outs_0_valid : std_logic;
  signal fork44_outs_0_ready : std_logic;
  signal fork44_outs_1 : std_logic_vector(31 downto 0);
  signal fork44_outs_1_valid : std_logic;
  signal fork44_outs_1_ready : std_logic;
  signal control_merge7_outs_valid : std_logic;
  signal control_merge7_outs_ready : std_logic;
  signal control_merge7_index : std_logic_vector(0 downto 0);
  signal control_merge7_index_valid : std_logic;
  signal control_merge7_index_ready : std_logic;
  signal fork45_outs_0 : std_logic_vector(0 downto 0);
  signal fork45_outs_0_valid : std_logic;
  signal fork45_outs_0_ready : std_logic;
  signal fork45_outs_1 : std_logic_vector(0 downto 0);
  signal fork45_outs_1_valid : std_logic;
  signal fork45_outs_1_ready : std_logic;
  signal fork45_outs_2 : std_logic_vector(0 downto 0);
  signal fork45_outs_2_valid : std_logic;
  signal fork45_outs_2_ready : std_logic;
  signal buffer100_outs_valid : std_logic;
  signal buffer100_outs_ready : std_logic;
  signal fork46_outs_0_valid : std_logic;
  signal fork46_outs_0_ready : std_logic;
  signal fork46_outs_1_valid : std_logic;
  signal fork46_outs_1_ready : std_logic;
  signal constant65_outs : std_logic_vector(1 downto 0);
  signal constant65_outs_valid : std_logic;
  signal constant65_outs_ready : std_logic;
  signal extsi22_outs : std_logic_vector(31 downto 0);
  signal extsi22_outs_valid : std_logic;
  signal extsi22_outs_ready : std_logic;
  signal source11_outs_valid : std_logic;
  signal source11_outs_ready : std_logic;
  signal constant66_outs : std_logic_vector(4 downto 0);
  signal constant66_outs_valid : std_logic;
  signal constant66_outs_ready : std_logic;
  signal extsi78_outs : std_logic_vector(5 downto 0);
  signal extsi78_outs_valid : std_logic;
  signal extsi78_outs_ready : std_logic;
  signal source12_outs_valid : std_logic;
  signal source12_outs_ready : std_logic;
  signal constant67_outs : std_logic_vector(1 downto 0);
  signal constant67_outs_valid : std_logic;
  signal constant67_outs_ready : std_logic;
  signal fork47_outs_0 : std_logic_vector(1 downto 0);
  signal fork47_outs_0_valid : std_logic;
  signal fork47_outs_0_ready : std_logic;
  signal fork47_outs_1 : std_logic_vector(1 downto 0);
  signal fork47_outs_1_valid : std_logic;
  signal fork47_outs_1_ready : std_logic;
  signal extsi79_outs : std_logic_vector(5 downto 0);
  signal extsi79_outs_valid : std_logic;
  signal extsi79_outs_ready : std_logic;
  signal extsi24_outs : std_logic_vector(31 downto 0);
  signal extsi24_outs_valid : std_logic;
  signal extsi24_outs_ready : std_logic;
  signal fork48_outs_0 : std_logic_vector(31 downto 0);
  signal fork48_outs_0_valid : std_logic;
  signal fork48_outs_0_ready : std_logic;
  signal fork48_outs_1 : std_logic_vector(31 downto 0);
  signal fork48_outs_1_valid : std_logic;
  signal fork48_outs_1_ready : std_logic;
  signal fork48_outs_2 : std_logic_vector(31 downto 0);
  signal fork48_outs_2_valid : std_logic;
  signal fork48_outs_2_ready : std_logic;
  signal fork48_outs_3 : std_logic_vector(31 downto 0);
  signal fork48_outs_3_valid : std_logic;
  signal fork48_outs_3_ready : std_logic;
  signal source13_outs_valid : std_logic;
  signal source13_outs_ready : std_logic;
  signal constant68_outs : std_logic_vector(2 downto 0);
  signal constant68_outs_valid : std_logic;
  signal constant68_outs_ready : std_logic;
  signal extsi25_outs : std_logic_vector(31 downto 0);
  signal extsi25_outs_valid : std_logic;
  signal extsi25_outs_ready : std_logic;
  signal fork49_outs_0 : std_logic_vector(31 downto 0);
  signal fork49_outs_0_valid : std_logic;
  signal fork49_outs_0_ready : std_logic;
  signal fork49_outs_1 : std_logic_vector(31 downto 0);
  signal fork49_outs_1_valid : std_logic;
  signal fork49_outs_1_ready : std_logic;
  signal fork49_outs_2 : std_logic_vector(31 downto 0);
  signal fork49_outs_2_valid : std_logic;
  signal fork49_outs_2_ready : std_logic;
  signal fork49_outs_3 : std_logic_vector(31 downto 0);
  signal fork49_outs_3_valid : std_logic;
  signal fork49_outs_3_ready : std_logic;
  signal shli12_result : std_logic_vector(31 downto 0);
  signal shli12_result_valid : std_logic;
  signal shli12_result_ready : std_logic;
  signal buffer103_outs : std_logic_vector(31 downto 0);
  signal buffer103_outs_valid : std_logic;
  signal buffer103_outs_ready : std_logic;
  signal buffer101_outs : std_logic_vector(31 downto 0);
  signal buffer101_outs_valid : std_logic;
  signal buffer101_outs_ready : std_logic;
  signal trunci13_outs : std_logic_vector(6 downto 0);
  signal trunci13_outs_valid : std_logic;
  signal trunci13_outs_ready : std_logic;
  signal shli13_result : std_logic_vector(31 downto 0);
  signal shli13_result_valid : std_logic;
  signal shli13_result_ready : std_logic;
  signal buffer105_outs : std_logic_vector(31 downto 0);
  signal buffer105_outs_valid : std_logic;
  signal buffer105_outs_ready : std_logic;
  signal buffer102_outs : std_logic_vector(31 downto 0);
  signal buffer102_outs_valid : std_logic;
  signal buffer102_outs_ready : std_logic;
  signal trunci14_outs : std_logic_vector(6 downto 0);
  signal trunci14_outs_valid : std_logic;
  signal trunci14_outs_ready : std_logic;
  signal addi33_result : std_logic_vector(6 downto 0);
  signal addi33_result_valid : std_logic;
  signal addi33_result_ready : std_logic;
  signal buffer104_outs : std_logic_vector(6 downto 0);
  signal buffer104_outs_valid : std_logic;
  signal buffer104_outs_ready : std_logic;
  signal addi9_result : std_logic_vector(6 downto 0);
  signal addi9_result_valid : std_logic;
  signal addi9_result_ready : std_logic;
  signal load3_addrOut : std_logic_vector(6 downto 0);
  signal load3_addrOut_valid : std_logic;
  signal load3_addrOut_ready : std_logic;
  signal load3_dataOut : std_logic_vector(31 downto 0);
  signal load3_dataOut_valid : std_logic;
  signal load3_dataOut_ready : std_logic;
  signal shli14_result : std_logic_vector(31 downto 0);
  signal shli14_result_valid : std_logic;
  signal shli14_result_ready : std_logic;
  signal buffer107_outs : std_logic_vector(31 downto 0);
  signal buffer107_outs_valid : std_logic;
  signal buffer107_outs_ready : std_logic;
  signal buffer106_outs : std_logic_vector(31 downto 0);
  signal buffer106_outs_valid : std_logic;
  signal buffer106_outs_ready : std_logic;
  signal trunci15_outs : std_logic_vector(6 downto 0);
  signal trunci15_outs_valid : std_logic;
  signal trunci15_outs_ready : std_logic;
  signal shli15_result : std_logic_vector(31 downto 0);
  signal shli15_result_valid : std_logic;
  signal shli15_result_ready : std_logic;
  signal buffer109_outs : std_logic_vector(31 downto 0);
  signal buffer109_outs_valid : std_logic;
  signal buffer109_outs_ready : std_logic;
  signal buffer108_outs : std_logic_vector(31 downto 0);
  signal buffer108_outs_valid : std_logic;
  signal buffer108_outs_ready : std_logic;
  signal trunci16_outs : std_logic_vector(6 downto 0);
  signal trunci16_outs_valid : std_logic;
  signal trunci16_outs_ready : std_logic;
  signal addi34_result : std_logic_vector(6 downto 0);
  signal addi34_result_valid : std_logic;
  signal addi34_result_ready : std_logic;
  signal buffer114_outs : std_logic_vector(6 downto 0);
  signal buffer114_outs_valid : std_logic;
  signal buffer114_outs_ready : std_logic;
  signal addi10_result : std_logic_vector(6 downto 0);
  signal addi10_result_valid : std_logic;
  signal addi10_result_ready : std_logic;
  signal load4_addrOut : std_logic_vector(6 downto 0);
  signal load4_addrOut_valid : std_logic;
  signal load4_addrOut_ready : std_logic;
  signal load4_dataOut : std_logic_vector(31 downto 0);
  signal load4_dataOut_valid : std_logic;
  signal load4_dataOut_ready : std_logic;
  signal muli1_result : std_logic_vector(31 downto 0);
  signal muli1_result_valid : std_logic;
  signal muli1_result_ready : std_logic;
  signal shli16_result : std_logic_vector(31 downto 0);
  signal shli16_result_valid : std_logic;
  signal shli16_result_ready : std_logic;
  signal buffer110_outs : std_logic_vector(31 downto 0);
  signal buffer110_outs_valid : std_logic;
  signal buffer110_outs_ready : std_logic;
  signal buffer111_outs : std_logic_vector(31 downto 0);
  signal buffer111_outs_valid : std_logic;
  signal buffer111_outs_ready : std_logic;
  signal shli17_result : std_logic_vector(31 downto 0);
  signal shli17_result_valid : std_logic;
  signal shli17_result_ready : std_logic;
  signal buffer112_outs : std_logic_vector(31 downto 0);
  signal buffer112_outs_valid : std_logic;
  signal buffer112_outs_ready : std_logic;
  signal buffer113_outs : std_logic_vector(31 downto 0);
  signal buffer113_outs_valid : std_logic;
  signal buffer113_outs_ready : std_logic;
  signal buffer119_outs : std_logic_vector(31 downto 0);
  signal buffer119_outs_valid : std_logic;
  signal buffer119_outs_ready : std_logic;
  signal buffer120_outs : std_logic_vector(31 downto 0);
  signal buffer120_outs_valid : std_logic;
  signal buffer120_outs_ready : std_logic;
  signal addi35_result : std_logic_vector(31 downto 0);
  signal addi35_result_valid : std_logic;
  signal addi35_result_ready : std_logic;
  signal buffer122_outs : std_logic_vector(31 downto 0);
  signal buffer122_outs_valid : std_logic;
  signal buffer122_outs_ready : std_logic;
  signal addi11_result : std_logic_vector(31 downto 0);
  signal addi11_result_valid : std_logic;
  signal addi11_result_ready : std_logic;
  signal buffer91_outs_valid : std_logic;
  signal buffer91_outs_ready : std_logic;
  signal gate2_outs : std_logic_vector(31 downto 0);
  signal gate2_outs_valid : std_logic;
  signal gate2_outs_ready : std_logic;
  signal trunci17_outs : std_logic_vector(6 downto 0);
  signal trunci17_outs_valid : std_logic;
  signal trunci17_outs_ready : std_logic;
  signal load5_addrOut : std_logic_vector(6 downto 0);
  signal load5_addrOut_valid : std_logic;
  signal load5_addrOut_ready : std_logic;
  signal load5_dataOut : std_logic_vector(31 downto 0);
  signal load5_dataOut_valid : std_logic;
  signal load5_dataOut_ready : std_logic;
  signal addi1_result : std_logic_vector(31 downto 0);
  signal addi1_result_valid : std_logic;
  signal addi1_result_ready : std_logic;
  signal shli18_result : std_logic_vector(31 downto 0);
  signal shli18_result_valid : std_logic;
  signal shli18_result_ready : std_logic;
  signal buffer115_outs : std_logic_vector(31 downto 0);
  signal buffer115_outs_valid : std_logic;
  signal buffer115_outs_ready : std_logic;
  signal buffer116_outs : std_logic_vector(31 downto 0);
  signal buffer116_outs_valid : std_logic;
  signal buffer116_outs_ready : std_logic;
  signal shli19_result : std_logic_vector(31 downto 0);
  signal shli19_result_valid : std_logic;
  signal shli19_result_ready : std_logic;
  signal buffer117_outs : std_logic_vector(31 downto 0);
  signal buffer117_outs_valid : std_logic;
  signal buffer117_outs_ready : std_logic;
  signal buffer118_outs : std_logic_vector(31 downto 0);
  signal buffer118_outs_valid : std_logic;
  signal buffer118_outs_ready : std_logic;
  signal buffer123_outs : std_logic_vector(31 downto 0);
  signal buffer123_outs_valid : std_logic;
  signal buffer123_outs_ready : std_logic;
  signal buffer124_outs : std_logic_vector(31 downto 0);
  signal buffer124_outs_valid : std_logic;
  signal buffer124_outs_ready : std_logic;
  signal addi36_result : std_logic_vector(31 downto 0);
  signal addi36_result_valid : std_logic;
  signal addi36_result_ready : std_logic;
  signal buffer125_outs : std_logic_vector(31 downto 0);
  signal buffer125_outs_valid : std_logic;
  signal buffer125_outs_ready : std_logic;
  signal addi12_result : std_logic_vector(31 downto 0);
  signal addi12_result_valid : std_logic;
  signal addi12_result_ready : std_logic;
  signal buffer3_outs_valid : std_logic;
  signal buffer3_outs_ready : std_logic;
  signal gate3_outs : std_logic_vector(31 downto 0);
  signal gate3_outs_valid : std_logic;
  signal gate3_outs_ready : std_logic;
  signal trunci18_outs : std_logic_vector(6 downto 0);
  signal trunci18_outs_valid : std_logic;
  signal trunci18_outs_ready : std_logic;
  signal store3_addrOut : std_logic_vector(6 downto 0);
  signal store3_addrOut_valid : std_logic;
  signal store3_addrOut_ready : std_logic;
  signal store3_dataToMem : std_logic_vector(31 downto 0);
  signal store3_dataToMem_valid : std_logic;
  signal store3_dataToMem_ready : std_logic;
  signal store3_doneOut_valid : std_logic;
  signal store3_doneOut_ready : std_logic;
  signal addi21_result : std_logic_vector(5 downto 0);
  signal addi21_result_valid : std_logic;
  signal addi21_result_ready : std_logic;
  signal fork50_outs_0 : std_logic_vector(5 downto 0);
  signal fork50_outs_0_valid : std_logic;
  signal fork50_outs_0_ready : std_logic;
  signal fork50_outs_1 : std_logic_vector(5 downto 0);
  signal fork50_outs_1_valid : std_logic;
  signal fork50_outs_1_ready : std_logic;
  signal trunci19_outs : std_logic_vector(4 downto 0);
  signal trunci19_outs_valid : std_logic;
  signal trunci19_outs_ready : std_logic;
  signal buffer131_outs : std_logic_vector(5 downto 0);
  signal buffer131_outs_valid : std_logic;
  signal buffer131_outs_ready : std_logic;
  signal cmpi3_result : std_logic_vector(0 downto 0);
  signal cmpi3_result_valid : std_logic;
  signal cmpi3_result_ready : std_logic;
  signal buffer121_outs : std_logic_vector(5 downto 0);
  signal buffer121_outs_valid : std_logic;
  signal buffer121_outs_ready : std_logic;
  signal buffer130_outs : std_logic_vector(0 downto 0);
  signal buffer130_outs_valid : std_logic;
  signal buffer130_outs_ready : std_logic;
  signal fork51_outs_0 : std_logic_vector(0 downto 0);
  signal fork51_outs_0_valid : std_logic;
  signal fork51_outs_0_ready : std_logic;
  signal fork51_outs_1 : std_logic_vector(0 downto 0);
  signal fork51_outs_1_valid : std_logic;
  signal fork51_outs_1_ready : std_logic;
  signal fork51_outs_2 : std_logic_vector(0 downto 0);
  signal fork51_outs_2_valid : std_logic;
  signal fork51_outs_2_ready : std_logic;
  signal fork51_outs_3 : std_logic_vector(0 downto 0);
  signal fork51_outs_3_valid : std_logic;
  signal fork51_outs_3_ready : std_logic;
  signal fork51_outs_4 : std_logic_vector(0 downto 0);
  signal fork51_outs_4_valid : std_logic;
  signal fork51_outs_4_ready : std_logic;
  signal fork51_outs_5 : std_logic_vector(0 downto 0);
  signal fork51_outs_5_valid : std_logic;
  signal fork51_outs_5_ready : std_logic;
  signal fork51_outs_6 : std_logic_vector(0 downto 0);
  signal fork51_outs_6_valid : std_logic;
  signal fork51_outs_6_ready : std_logic;
  signal cond_br19_trueOut : std_logic_vector(4 downto 0);
  signal cond_br19_trueOut_valid : std_logic;
  signal cond_br19_trueOut_ready : std_logic;
  signal cond_br19_falseOut : std_logic_vector(4 downto 0);
  signal cond_br19_falseOut_valid : std_logic;
  signal cond_br19_falseOut_ready : std_logic;
  signal cond_br20_trueOut : std_logic_vector(4 downto 0);
  signal cond_br20_trueOut_valid : std_logic;
  signal cond_br20_trueOut_ready : std_logic;
  signal cond_br20_falseOut : std_logic_vector(4 downto 0);
  signal cond_br20_falseOut_valid : std_logic;
  signal cond_br20_falseOut_ready : std_logic;
  signal cond_br21_trueOut : std_logic_vector(4 downto 0);
  signal cond_br21_trueOut_valid : std_logic;
  signal cond_br21_trueOut_ready : std_logic;
  signal cond_br21_falseOut : std_logic_vector(4 downto 0);
  signal cond_br21_falseOut_valid : std_logic;
  signal cond_br21_falseOut_ready : std_logic;
  signal cond_br22_trueOut_valid : std_logic;
  signal cond_br22_trueOut_ready : std_logic;
  signal cond_br22_falseOut_valid : std_logic;
  signal cond_br22_falseOut_ready : std_logic;
  signal buffer127_outs : std_logic_vector(0 downto 0);
  signal buffer127_outs_valid : std_logic;
  signal buffer127_outs_ready : std_logic;
  signal cond_br124_trueOut_valid : std_logic;
  signal cond_br124_trueOut_ready : std_logic;
  signal cond_br124_falseOut_valid : std_logic;
  signal cond_br124_falseOut_ready : std_logic;
  signal buffer128_outs : std_logic_vector(0 downto 0);
  signal buffer128_outs_valid : std_logic;
  signal buffer128_outs_ready : std_logic;
  signal cond_br125_trueOut_valid : std_logic;
  signal cond_br125_trueOut_ready : std_logic;
  signal cond_br125_falseOut_valid : std_logic;
  signal cond_br125_falseOut_ready : std_logic;
  signal buffer129_outs : std_logic_vector(0 downto 0);
  signal buffer129_outs_valid : std_logic;
  signal buffer129_outs_ready : std_logic;
  signal extsi80_outs : std_logic_vector(5 downto 0);
  signal extsi80_outs_valid : std_logic;
  signal extsi80_outs_ready : std_logic;
  signal source14_outs_valid : std_logic;
  signal source14_outs_ready : std_logic;
  signal constant69_outs : std_logic_vector(4 downto 0);
  signal constant69_outs_valid : std_logic;
  signal constant69_outs_ready : std_logic;
  signal extsi81_outs : std_logic_vector(5 downto 0);
  signal extsi81_outs_valid : std_logic;
  signal extsi81_outs_ready : std_logic;
  signal source15_outs_valid : std_logic;
  signal source15_outs_ready : std_logic;
  signal constant70_outs : std_logic_vector(1 downto 0);
  signal constant70_outs_valid : std_logic;
  signal constant70_outs_ready : std_logic;
  signal extsi82_outs : std_logic_vector(5 downto 0);
  signal extsi82_outs_valid : std_logic;
  signal extsi82_outs_ready : std_logic;
  signal addi22_result : std_logic_vector(5 downto 0);
  signal addi22_result_valid : std_logic;
  signal addi22_result_ready : std_logic;
  signal buffer132_outs : std_logic_vector(5 downto 0);
  signal buffer132_outs_valid : std_logic;
  signal buffer132_outs_ready : std_logic;
  signal fork52_outs_0 : std_logic_vector(5 downto 0);
  signal fork52_outs_0_valid : std_logic;
  signal fork52_outs_0_ready : std_logic;
  signal fork52_outs_1 : std_logic_vector(5 downto 0);
  signal fork52_outs_1_valid : std_logic;
  signal fork52_outs_1_ready : std_logic;
  signal trunci20_outs : std_logic_vector(4 downto 0);
  signal trunci20_outs_valid : std_logic;
  signal trunci20_outs_ready : std_logic;
  signal cmpi4_result : std_logic_vector(0 downto 0);
  signal cmpi4_result_valid : std_logic;
  signal cmpi4_result_ready : std_logic;
  signal buffer133_outs : std_logic_vector(0 downto 0);
  signal buffer133_outs_valid : std_logic;
  signal buffer133_outs_ready : std_logic;
  signal fork53_outs_0 : std_logic_vector(0 downto 0);
  signal fork53_outs_0_valid : std_logic;
  signal fork53_outs_0_ready : std_logic;
  signal fork53_outs_1 : std_logic_vector(0 downto 0);
  signal fork53_outs_1_valid : std_logic;
  signal fork53_outs_1_ready : std_logic;
  signal fork53_outs_2 : std_logic_vector(0 downto 0);
  signal fork53_outs_2_valid : std_logic;
  signal fork53_outs_2_ready : std_logic;
  signal fork53_outs_3 : std_logic_vector(0 downto 0);
  signal fork53_outs_3_valid : std_logic;
  signal fork53_outs_3_ready : std_logic;
  signal fork53_outs_4 : std_logic_vector(0 downto 0);
  signal fork53_outs_4_valid : std_logic;
  signal fork53_outs_4_ready : std_logic;
  signal fork53_outs_5 : std_logic_vector(0 downto 0);
  signal fork53_outs_5_valid : std_logic;
  signal fork53_outs_5_ready : std_logic;
  signal cond_br23_trueOut : std_logic_vector(4 downto 0);
  signal cond_br23_trueOut_valid : std_logic;
  signal cond_br23_trueOut_ready : std_logic;
  signal cond_br23_falseOut : std_logic_vector(4 downto 0);
  signal cond_br23_falseOut_valid : std_logic;
  signal cond_br23_falseOut_ready : std_logic;
  signal cond_br24_trueOut : std_logic_vector(4 downto 0);
  signal cond_br24_trueOut_valid : std_logic;
  signal cond_br24_trueOut_ready : std_logic;
  signal cond_br24_falseOut : std_logic_vector(4 downto 0);
  signal cond_br24_falseOut_valid : std_logic;
  signal cond_br24_falseOut_ready : std_logic;
  signal cond_br25_trueOut_valid : std_logic;
  signal cond_br25_trueOut_ready : std_logic;
  signal cond_br25_falseOut_valid : std_logic;
  signal cond_br25_falseOut_ready : std_logic;
  signal buffer134_outs : std_logic_vector(0 downto 0);
  signal buffer134_outs_valid : std_logic;
  signal buffer134_outs_ready : std_logic;
  signal cond_br126_trueOut_valid : std_logic;
  signal cond_br126_trueOut_ready : std_logic;
  signal cond_br126_falseOut_valid : std_logic;
  signal cond_br126_falseOut_ready : std_logic;
  signal cond_br127_trueOut_valid : std_logic;
  signal cond_br127_trueOut_ready : std_logic;
  signal cond_br127_falseOut_valid : std_logic;
  signal cond_br127_falseOut_ready : std_logic;
  signal buffer136_outs : std_logic_vector(0 downto 0);
  signal buffer136_outs_valid : std_logic;
  signal buffer136_outs_ready : std_logic;
  signal buffer135_outs : std_logic_vector(4 downto 0);
  signal buffer135_outs_valid : std_logic;
  signal buffer135_outs_ready : std_logic;
  signal extsi83_outs : std_logic_vector(5 downto 0);
  signal extsi83_outs_valid : std_logic;
  signal extsi83_outs_ready : std_logic;
  signal fork54_outs_0_valid : std_logic;
  signal fork54_outs_0_ready : std_logic;
  signal fork54_outs_1_valid : std_logic;
  signal fork54_outs_1_ready : std_logic;
  signal constant71_outs : std_logic_vector(0 downto 0);
  signal constant71_outs_valid : std_logic;
  signal constant71_outs_ready : std_logic;
  signal source16_outs_valid : std_logic;
  signal source16_outs_ready : std_logic;
  signal constant72_outs : std_logic_vector(4 downto 0);
  signal constant72_outs_valid : std_logic;
  signal constant72_outs_ready : std_logic;
  signal extsi84_outs : std_logic_vector(5 downto 0);
  signal extsi84_outs_valid : std_logic;
  signal extsi84_outs_ready : std_logic;
  signal source17_outs_valid : std_logic;
  signal source17_outs_ready : std_logic;
  signal constant73_outs : std_logic_vector(1 downto 0);
  signal constant73_outs_valid : std_logic;
  signal constant73_outs_ready : std_logic;
  signal extsi85_outs : std_logic_vector(5 downto 0);
  signal extsi85_outs_valid : std_logic;
  signal extsi85_outs_ready : std_logic;
  signal addi23_result : std_logic_vector(5 downto 0);
  signal addi23_result_valid : std_logic;
  signal addi23_result_ready : std_logic;
  signal buffer137_outs : std_logic_vector(5 downto 0);
  signal buffer137_outs_valid : std_logic;
  signal buffer137_outs_ready : std_logic;
  signal fork55_outs_0 : std_logic_vector(5 downto 0);
  signal fork55_outs_0_valid : std_logic;
  signal fork55_outs_0_ready : std_logic;
  signal fork55_outs_1 : std_logic_vector(5 downto 0);
  signal fork55_outs_1_valid : std_logic;
  signal fork55_outs_1_ready : std_logic;
  signal trunci21_outs : std_logic_vector(4 downto 0);
  signal trunci21_outs_valid : std_logic;
  signal trunci21_outs_ready : std_logic;
  signal cmpi5_result : std_logic_vector(0 downto 0);
  signal cmpi5_result_valid : std_logic;
  signal cmpi5_result_ready : std_logic;
  signal buffer138_outs : std_logic_vector(0 downto 0);
  signal buffer138_outs_valid : std_logic;
  signal buffer138_outs_ready : std_logic;
  signal fork56_outs_0 : std_logic_vector(0 downto 0);
  signal fork56_outs_0_valid : std_logic;
  signal fork56_outs_0_ready : std_logic;
  signal fork56_outs_1 : std_logic_vector(0 downto 0);
  signal fork56_outs_1_valid : std_logic;
  signal fork56_outs_1_ready : std_logic;
  signal fork56_outs_2 : std_logic_vector(0 downto 0);
  signal fork56_outs_2_valid : std_logic;
  signal fork56_outs_2_ready : std_logic;
  signal fork56_outs_3 : std_logic_vector(0 downto 0);
  signal fork56_outs_3_valid : std_logic;
  signal fork56_outs_3_ready : std_logic;
  signal fork56_outs_4 : std_logic_vector(0 downto 0);
  signal fork56_outs_4_valid : std_logic;
  signal fork56_outs_4_ready : std_logic;
  signal fork56_outs_5 : std_logic_vector(0 downto 0);
  signal fork56_outs_5_valid : std_logic;
  signal fork56_outs_5_ready : std_logic;
  signal cond_br26_trueOut : std_logic_vector(4 downto 0);
  signal cond_br26_trueOut_valid : std_logic;
  signal cond_br26_trueOut_ready : std_logic;
  signal cond_br26_falseOut : std_logic_vector(4 downto 0);
  signal cond_br26_falseOut_valid : std_logic;
  signal cond_br26_falseOut_ready : std_logic;
  signal cond_br27_trueOut_valid : std_logic;
  signal cond_br27_trueOut_ready : std_logic;
  signal cond_br27_falseOut_valid : std_logic;
  signal cond_br27_falseOut_ready : std_logic;
  signal cond_br28_trueOut : std_logic_vector(0 downto 0);
  signal cond_br28_trueOut_valid : std_logic;
  signal cond_br28_trueOut_ready : std_logic;
  signal cond_br28_falseOut : std_logic_vector(0 downto 0);
  signal cond_br28_falseOut_valid : std_logic;
  signal cond_br28_falseOut_ready : std_logic;
  signal extsi47_outs : std_logic_vector(4 downto 0);
  signal extsi47_outs_valid : std_logic;
  signal extsi47_outs_ready : std_logic;
  signal init28_outs : std_logic_vector(0 downto 0);
  signal init28_outs_valid : std_logic;
  signal init28_outs_ready : std_logic;
  signal fork57_outs_0 : std_logic_vector(0 downto 0);
  signal fork57_outs_0_valid : std_logic;
  signal fork57_outs_0_ready : std_logic;
  signal fork57_outs_1 : std_logic_vector(0 downto 0);
  signal fork57_outs_1_valid : std_logic;
  signal fork57_outs_1_ready : std_logic;
  signal fork57_outs_2 : std_logic_vector(0 downto 0);
  signal fork57_outs_2_valid : std_logic;
  signal fork57_outs_2_ready : std_logic;
  signal fork57_outs_3 : std_logic_vector(0 downto 0);
  signal fork57_outs_3_valid : std_logic;
  signal fork57_outs_3_ready : std_logic;
  signal fork57_outs_4 : std_logic_vector(0 downto 0);
  signal fork57_outs_4_valid : std_logic;
  signal fork57_outs_4_ready : std_logic;
  signal mux46_outs_valid : std_logic;
  signal mux46_outs_ready : std_logic;
  signal buffer143_outs : std_logic_vector(0 downto 0);
  signal buffer143_outs_valid : std_logic;
  signal buffer143_outs_ready : std_logic;
  signal buffer139_outs_valid : std_logic;
  signal buffer139_outs_ready : std_logic;
  signal buffer140_outs_valid : std_logic;
  signal buffer140_outs_ready : std_logic;
  signal fork58_outs_0_valid : std_logic;
  signal fork58_outs_0_ready : std_logic;
  signal fork58_outs_1_valid : std_logic;
  signal fork58_outs_1_ready : std_logic;
  signal mux47_outs_valid : std_logic;
  signal mux47_outs_ready : std_logic;
  signal buffer144_outs : std_logic_vector(0 downto 0);
  signal buffer144_outs_valid : std_logic;
  signal buffer144_outs_ready : std_logic;
  signal buffer141_outs_valid : std_logic;
  signal buffer141_outs_ready : std_logic;
  signal buffer142_outs_valid : std_logic;
  signal buffer142_outs_ready : std_logic;
  signal fork59_outs_0_valid : std_logic;
  signal fork59_outs_0_ready : std_logic;
  signal fork59_outs_1_valid : std_logic;
  signal fork59_outs_1_ready : std_logic;
  signal buffer245_outs_valid : std_logic;
  signal buffer245_outs_ready : std_logic;
  signal mux48_outs_valid : std_logic;
  signal mux48_outs_ready : std_logic;
  signal buffer145_outs : std_logic_vector(0 downto 0);
  signal buffer145_outs_valid : std_logic;
  signal buffer145_outs_ready : std_logic;
  signal buffer146_outs_valid : std_logic;
  signal buffer146_outs_ready : std_logic;
  signal fork60_outs_0_valid : std_logic;
  signal fork60_outs_0_ready : std_logic;
  signal fork60_outs_1_valid : std_logic;
  signal fork60_outs_1_ready : std_logic;
  signal mux49_outs_valid : std_logic;
  signal mux49_outs_ready : std_logic;
  signal buffer147_outs_valid : std_logic;
  signal buffer147_outs_ready : std_logic;
  signal buffer148_outs_valid : std_logic;
  signal buffer148_outs_ready : std_logic;
  signal fork61_outs_0_valid : std_logic;
  signal fork61_outs_0_ready : std_logic;
  signal fork61_outs_1_valid : std_logic;
  signal fork61_outs_1_ready : std_logic;
  signal mux51_outs_valid : std_logic;
  signal mux51_outs_ready : std_logic;
  signal mux12_outs : std_logic_vector(4 downto 0);
  signal mux12_outs_valid : std_logic;
  signal mux12_outs_ready : std_logic;
  signal control_merge10_outs_valid : std_logic;
  signal control_merge10_outs_ready : std_logic;
  signal control_merge10_index : std_logic_vector(0 downto 0);
  signal control_merge10_index_valid : std_logic;
  signal control_merge10_index_ready : std_logic;
  signal fork62_outs_0_valid : std_logic;
  signal fork62_outs_0_ready : std_logic;
  signal fork62_outs_1_valid : std_logic;
  signal fork62_outs_1_ready : std_logic;
  signal constant74_outs : std_logic_vector(0 downto 0);
  signal constant74_outs_valid : std_logic;
  signal constant74_outs_ready : std_logic;
  signal extsi46_outs : std_logic_vector(4 downto 0);
  signal extsi46_outs_valid : std_logic;
  signal extsi46_outs_ready : std_logic;
  signal buffer151_outs : std_logic_vector(4 downto 0);
  signal buffer151_outs_valid : std_logic;
  signal buffer151_outs_ready : std_logic;
  signal init35_outs : std_logic_vector(0 downto 0);
  signal init35_outs_valid : std_logic;
  signal init35_outs_ready : std_logic;
  signal fork63_outs_0 : std_logic_vector(0 downto 0);
  signal fork63_outs_0_valid : std_logic;
  signal fork63_outs_0_ready : std_logic;
  signal fork63_outs_1 : std_logic_vector(0 downto 0);
  signal fork63_outs_1_valid : std_logic;
  signal fork63_outs_1_ready : std_logic;
  signal fork63_outs_2 : std_logic_vector(0 downto 0);
  signal fork63_outs_2_valid : std_logic;
  signal fork63_outs_2_ready : std_logic;
  signal fork63_outs_3 : std_logic_vector(0 downto 0);
  signal fork63_outs_3_valid : std_logic;
  signal fork63_outs_3_ready : std_logic;
  signal fork63_outs_4 : std_logic_vector(0 downto 0);
  signal fork63_outs_4_valid : std_logic;
  signal fork63_outs_4_ready : std_logic;
  signal mux53_outs_valid : std_logic;
  signal mux53_outs_ready : std_logic;
  signal buffer152_outs_valid : std_logic;
  signal buffer152_outs_ready : std_logic;
  signal buffer154_outs_valid : std_logic;
  signal buffer154_outs_ready : std_logic;
  signal fork64_outs_0_valid : std_logic;
  signal fork64_outs_0_ready : std_logic;
  signal fork64_outs_1_valid : std_logic;
  signal fork64_outs_1_ready : std_logic;
  signal buffer242_outs_valid : std_logic;
  signal buffer242_outs_ready : std_logic;
  signal mux54_outs_valid : std_logic;
  signal mux54_outs_ready : std_logic;
  signal buffer155_outs_valid : std_logic;
  signal buffer155_outs_ready : std_logic;
  signal fork65_outs_0_valid : std_logic;
  signal fork65_outs_0_ready : std_logic;
  signal fork65_outs_1_valid : std_logic;
  signal fork65_outs_1_ready : std_logic;
  signal mux55_outs_valid : std_logic;
  signal mux55_outs_ready : std_logic;
  signal buffer156_outs_valid : std_logic;
  signal buffer156_outs_ready : std_logic;
  signal buffer157_outs_valid : std_logic;
  signal buffer157_outs_ready : std_logic;
  signal fork66_outs_0_valid : std_logic;
  signal fork66_outs_0_ready : std_logic;
  signal fork66_outs_1_valid : std_logic;
  signal fork66_outs_1_ready : std_logic;
  signal mux56_outs_valid : std_logic;
  signal mux56_outs_ready : std_logic;
  signal buffer158_outs_valid : std_logic;
  signal buffer158_outs_ready : std_logic;
  signal buffer159_outs_valid : std_logic;
  signal buffer159_outs_ready : std_logic;
  signal fork67_outs_0_valid : std_logic;
  signal fork67_outs_0_ready : std_logic;
  signal fork67_outs_1_valid : std_logic;
  signal fork67_outs_1_ready : std_logic;
  signal buffer149_outs_valid : std_logic;
  signal buffer149_outs_ready : std_logic;
  signal buffer150_outs_valid : std_logic;
  signal buffer150_outs_ready : std_logic;
  signal mux58_outs_valid : std_logic;
  signal mux58_outs_ready : std_logic;
  signal buffer153_outs : std_logic_vector(0 downto 0);
  signal buffer153_outs_valid : std_logic;
  signal buffer153_outs_ready : std_logic;
  signal mux13_outs : std_logic_vector(4 downto 0);
  signal mux13_outs_valid : std_logic;
  signal mux13_outs_ready : std_logic;
  signal buffer161_outs : std_logic_vector(4 downto 0);
  signal buffer161_outs_valid : std_logic;
  signal buffer161_outs_ready : std_logic;
  signal fork68_outs_0 : std_logic_vector(4 downto 0);
  signal fork68_outs_0_valid : std_logic;
  signal fork68_outs_0_ready : std_logic;
  signal fork68_outs_1 : std_logic_vector(4 downto 0);
  signal fork68_outs_1_valid : std_logic;
  signal fork68_outs_1_ready : std_logic;
  signal extsi86_outs : std_logic_vector(6 downto 0);
  signal extsi86_outs_valid : std_logic;
  signal extsi86_outs_ready : std_logic;
  signal mux14_outs : std_logic_vector(4 downto 0);
  signal mux14_outs_valid : std_logic;
  signal mux14_outs_ready : std_logic;
  signal buffer162_outs : std_logic_vector(4 downto 0);
  signal buffer162_outs_valid : std_logic;
  signal buffer162_outs_ready : std_logic;
  signal buffer163_outs : std_logic_vector(4 downto 0);
  signal buffer163_outs_valid : std_logic;
  signal buffer163_outs_ready : std_logic;
  signal fork69_outs_0 : std_logic_vector(4 downto 0);
  signal fork69_outs_0_valid : std_logic;
  signal fork69_outs_0_ready : std_logic;
  signal fork69_outs_1 : std_logic_vector(4 downto 0);
  signal fork69_outs_1_valid : std_logic;
  signal fork69_outs_1_ready : std_logic;
  signal extsi87_outs : std_logic_vector(31 downto 0);
  signal extsi87_outs_valid : std_logic;
  signal extsi87_outs_ready : std_logic;
  signal fork70_outs_0 : std_logic_vector(31 downto 0);
  signal fork70_outs_0_valid : std_logic;
  signal fork70_outs_0_ready : std_logic;
  signal fork70_outs_1 : std_logic_vector(31 downto 0);
  signal fork70_outs_1_valid : std_logic;
  signal fork70_outs_1_ready : std_logic;
  signal control_merge11_outs_valid : std_logic;
  signal control_merge11_outs_ready : std_logic;
  signal control_merge11_index : std_logic_vector(0 downto 0);
  signal control_merge11_index_valid : std_logic;
  signal control_merge11_index_ready : std_logic;
  signal fork71_outs_0 : std_logic_vector(0 downto 0);
  signal fork71_outs_0_valid : std_logic;
  signal fork71_outs_0_ready : std_logic;
  signal fork71_outs_1 : std_logic_vector(0 downto 0);
  signal fork71_outs_1_valid : std_logic;
  signal fork71_outs_1_ready : std_logic;
  signal fork72_outs_0_valid : std_logic;
  signal fork72_outs_0_ready : std_logic;
  signal fork72_outs_1_valid : std_logic;
  signal fork72_outs_1_ready : std_logic;
  signal fork72_outs_2_valid : std_logic;
  signal fork72_outs_2_ready : std_logic;
  signal constant75_outs : std_logic_vector(1 downto 0);
  signal constant75_outs_valid : std_logic;
  signal constant75_outs_ready : std_logic;
  signal extsi32_outs : std_logic_vector(31 downto 0);
  signal extsi32_outs_valid : std_logic;
  signal extsi32_outs_ready : std_logic;
  signal constant76_outs : std_logic_vector(0 downto 0);
  signal constant76_outs_valid : std_logic;
  signal constant76_outs_ready : std_logic;
  signal fork73_outs_0 : std_logic_vector(0 downto 0);
  signal fork73_outs_0_valid : std_logic;
  signal fork73_outs_0_ready : std_logic;
  signal fork73_outs_1 : std_logic_vector(0 downto 0);
  signal fork73_outs_1_valid : std_logic;
  signal fork73_outs_1_ready : std_logic;
  signal extsi34_outs : std_logic_vector(31 downto 0);
  signal extsi34_outs_valid : std_logic;
  signal extsi34_outs_ready : std_logic;
  signal source18_outs_valid : std_logic;
  signal source18_outs_ready : std_logic;
  signal constant77_outs : std_logic_vector(1 downto 0);
  signal constant77_outs_valid : std_logic;
  signal constant77_outs_ready : std_logic;
  signal extsi35_outs : std_logic_vector(31 downto 0);
  signal extsi35_outs_valid : std_logic;
  signal extsi35_outs_ready : std_logic;
  signal source19_outs_valid : std_logic;
  signal source19_outs_ready : std_logic;
  signal constant78_outs : std_logic_vector(2 downto 0);
  signal constant78_outs_valid : std_logic;
  signal constant78_outs_ready : std_logic;
  signal extsi36_outs : std_logic_vector(31 downto 0);
  signal extsi36_outs_valid : std_logic;
  signal extsi36_outs_ready : std_logic;
  signal shli20_result : std_logic_vector(31 downto 0);
  signal shli20_result_valid : std_logic;
  signal shli20_result_ready : std_logic;
  signal buffer170_outs : std_logic_vector(31 downto 0);
  signal buffer170_outs_valid : std_logic;
  signal buffer170_outs_ready : std_logic;
  signal trunci22_outs : std_logic_vector(6 downto 0);
  signal trunci22_outs_valid : std_logic;
  signal trunci22_outs_ready : std_logic;
  signal shli21_result : std_logic_vector(31 downto 0);
  signal shli21_result_valid : std_logic;
  signal shli21_result_ready : std_logic;
  signal buffer177_outs : std_logic_vector(31 downto 0);
  signal buffer177_outs_valid : std_logic;
  signal buffer177_outs_ready : std_logic;
  signal trunci23_outs : std_logic_vector(6 downto 0);
  signal trunci23_outs_valid : std_logic;
  signal trunci23_outs_ready : std_logic;
  signal addi37_result : std_logic_vector(6 downto 0);
  signal addi37_result_valid : std_logic;
  signal addi37_result_ready : std_logic;
  signal buffer178_outs : std_logic_vector(6 downto 0);
  signal buffer178_outs_valid : std_logic;
  signal buffer178_outs_ready : std_logic;
  signal addi13_result : std_logic_vector(6 downto 0);
  signal addi13_result_valid : std_logic;
  signal addi13_result_ready : std_logic;
  signal buffer4_outs_valid : std_logic;
  signal buffer4_outs_ready : std_logic;
  signal buffer179_outs : std_logic_vector(6 downto 0);
  signal buffer179_outs_valid : std_logic;
  signal buffer179_outs_ready : std_logic;
  signal store4_addrOut : std_logic_vector(6 downto 0);
  signal store4_addrOut_valid : std_logic;
  signal store4_addrOut_ready : std_logic;
  signal store4_dataToMem : std_logic_vector(31 downto 0);
  signal store4_dataToMem_valid : std_logic;
  signal store4_dataToMem_ready : std_logic;
  signal store4_doneOut_valid : std_logic;
  signal store4_doneOut_ready : std_logic;
  signal extsi45_outs : std_logic_vector(4 downto 0);
  signal extsi45_outs_valid : std_logic;
  signal extsi45_outs_ready : std_logic;
  signal buffer208_outs_valid : std_logic;
  signal buffer208_outs_ready : std_logic;
  signal cond_br128_trueOut_valid : std_logic;
  signal cond_br128_trueOut_ready : std_logic;
  signal cond_br128_falseOut_valid : std_logic;
  signal cond_br128_falseOut_ready : std_logic;
  signal buffer164_outs : std_logic_vector(0 downto 0);
  signal buffer164_outs_valid : std_logic;
  signal buffer164_outs_ready : std_logic;
  signal cond_br129_trueOut_valid : std_logic;
  signal cond_br129_trueOut_ready : std_logic;
  signal cond_br129_falseOut_valid : std_logic;
  signal cond_br129_falseOut_ready : std_logic;
  signal buffer165_outs : std_logic_vector(0 downto 0);
  signal buffer165_outs_valid : std_logic;
  signal buffer165_outs_ready : std_logic;
  signal cond_br130_trueOut_valid : std_logic;
  signal cond_br130_trueOut_ready : std_logic;
  signal cond_br130_falseOut_valid : std_logic;
  signal cond_br130_falseOut_ready : std_logic;
  signal buffer166_outs : std_logic_vector(0 downto 0);
  signal buffer166_outs_valid : std_logic;
  signal buffer166_outs_ready : std_logic;
  signal cond_br131_trueOut_valid : std_logic;
  signal cond_br131_trueOut_ready : std_logic;
  signal cond_br131_falseOut_valid : std_logic;
  signal cond_br131_falseOut_ready : std_logic;
  signal buffer167_outs : std_logic_vector(0 downto 0);
  signal buffer167_outs_valid : std_logic;
  signal buffer167_outs_ready : std_logic;
  signal cond_br132_trueOut_valid : std_logic;
  signal cond_br132_trueOut_ready : std_logic;
  signal cond_br132_falseOut_valid : std_logic;
  signal cond_br132_falseOut_ready : std_logic;
  signal buffer168_outs : std_logic_vector(0 downto 0);
  signal buffer168_outs_valid : std_logic;
  signal buffer168_outs_ready : std_logic;
  signal cond_br133_trueOut_valid : std_logic;
  signal cond_br133_trueOut_ready : std_logic;
  signal cond_br133_falseOut_valid : std_logic;
  signal cond_br133_falseOut_ready : std_logic;
  signal buffer169_outs : std_logic_vector(0 downto 0);
  signal buffer169_outs_valid : std_logic;
  signal buffer169_outs_ready : std_logic;
  signal init42_outs : std_logic_vector(0 downto 0);
  signal init42_outs_valid : std_logic;
  signal init42_outs_ready : std_logic;
  signal fork74_outs_0 : std_logic_vector(0 downto 0);
  signal fork74_outs_0_valid : std_logic;
  signal fork74_outs_0_ready : std_logic;
  signal fork74_outs_1 : std_logic_vector(0 downto 0);
  signal fork74_outs_1_valid : std_logic;
  signal fork74_outs_1_ready : std_logic;
  signal fork74_outs_2 : std_logic_vector(0 downto 0);
  signal fork74_outs_2_valid : std_logic;
  signal fork74_outs_2_ready : std_logic;
  signal fork74_outs_3 : std_logic_vector(0 downto 0);
  signal fork74_outs_3_valid : std_logic;
  signal fork74_outs_3_ready : std_logic;
  signal fork74_outs_4 : std_logic_vector(0 downto 0);
  signal fork74_outs_4_valid : std_logic;
  signal fork74_outs_4_ready : std_logic;
  signal fork74_outs_5 : std_logic_vector(0 downto 0);
  signal fork74_outs_5_valid : std_logic;
  signal fork74_outs_5_ready : std_logic;
  signal mux60_outs_valid : std_logic;
  signal mux60_outs_ready : std_logic;
  signal buffer171_outs : std_logic_vector(0 downto 0);
  signal buffer171_outs_valid : std_logic;
  signal buffer171_outs_ready : std_logic;
  signal buffer183_outs_valid : std_logic;
  signal buffer183_outs_ready : std_logic;
  signal buffer184_outs_valid : std_logic;
  signal buffer184_outs_ready : std_logic;
  signal fork75_outs_0_valid : std_logic;
  signal fork75_outs_0_ready : std_logic;
  signal fork75_outs_1_valid : std_logic;
  signal fork75_outs_1_ready : std_logic;
  signal fork75_outs_2_valid : std_logic;
  signal fork75_outs_2_ready : std_logic;
  signal buffer180_outs_valid : std_logic;
  signal buffer180_outs_ready : std_logic;
  signal mux62_outs_valid : std_logic;
  signal mux62_outs_ready : std_logic;
  signal buffer172_outs : std_logic_vector(0 downto 0);
  signal buffer172_outs_valid : std_logic;
  signal buffer172_outs_ready : std_logic;
  signal buffer186_outs_valid : std_logic;
  signal buffer186_outs_ready : std_logic;
  signal fork76_outs_0_valid : std_logic;
  signal fork76_outs_0_ready : std_logic;
  signal fork76_outs_1_valid : std_logic;
  signal fork76_outs_1_ready : std_logic;
  signal buffer182_outs_valid : std_logic;
  signal buffer182_outs_ready : std_logic;
  signal mux63_outs_valid : std_logic;
  signal mux63_outs_ready : std_logic;
  signal buffer173_outs : std_logic_vector(0 downto 0);
  signal buffer173_outs_valid : std_logic;
  signal buffer173_outs_ready : std_logic;
  signal buffer188_outs_valid : std_logic;
  signal buffer188_outs_ready : std_logic;
  signal fork77_outs_0_valid : std_logic;
  signal fork77_outs_0_ready : std_logic;
  signal fork77_outs_1_valid : std_logic;
  signal fork77_outs_1_ready : std_logic;
  signal mux64_outs_valid : std_logic;
  signal mux64_outs_ready : std_logic;
  signal buffer174_outs : std_logic_vector(0 downto 0);
  signal buffer174_outs_valid : std_logic;
  signal buffer174_outs_ready : std_logic;
  signal buffer191_outs_valid : std_logic;
  signal buffer191_outs_ready : std_logic;
  signal buffer193_outs_valid : std_logic;
  signal buffer193_outs_ready : std_logic;
  signal fork78_outs_0_valid : std_logic;
  signal fork78_outs_0_ready : std_logic;
  signal fork78_outs_1_valid : std_logic;
  signal fork78_outs_1_ready : std_logic;
  signal mux65_outs_valid : std_logic;
  signal mux65_outs_ready : std_logic;
  signal buffer175_outs : std_logic_vector(0 downto 0);
  signal buffer175_outs_valid : std_logic;
  signal buffer175_outs_ready : std_logic;
  signal buffer195_outs_valid : std_logic;
  signal buffer195_outs_ready : std_logic;
  signal fork79_outs_0_valid : std_logic;
  signal fork79_outs_0_ready : std_logic;
  signal fork79_outs_1_valid : std_logic;
  signal fork79_outs_1_ready : std_logic;
  signal buffer160_outs_valid : std_logic;
  signal buffer160_outs_ready : std_logic;
  signal mux66_outs_valid : std_logic;
  signal mux66_outs_ready : std_logic;
  signal buffer176_outs : std_logic_vector(0 downto 0);
  signal buffer176_outs_valid : std_logic;
  signal buffer176_outs_ready : std_logic;
  signal mux15_outs : std_logic_vector(4 downto 0);
  signal mux15_outs_valid : std_logic;
  signal mux15_outs_ready : std_logic;
  signal buffer215_outs : std_logic_vector(4 downto 0);
  signal buffer215_outs_valid : std_logic;
  signal buffer215_outs_ready : std_logic;
  signal buffer216_outs : std_logic_vector(4 downto 0);
  signal buffer216_outs_valid : std_logic;
  signal buffer216_outs_ready : std_logic;
  signal fork80_outs_0 : std_logic_vector(4 downto 0);
  signal fork80_outs_0_valid : std_logic;
  signal fork80_outs_0_ready : std_logic;
  signal fork80_outs_1 : std_logic_vector(4 downto 0);
  signal fork80_outs_1_valid : std_logic;
  signal fork80_outs_1_ready : std_logic;
  signal extsi88_outs : std_logic_vector(5 downto 0);
  signal extsi88_outs_valid : std_logic;
  signal extsi88_outs_ready : std_logic;
  signal extsi89_outs : std_logic_vector(31 downto 0);
  signal extsi89_outs_valid : std_logic;
  signal extsi89_outs_ready : std_logic;
  signal fork81_outs_0 : std_logic_vector(31 downto 0);
  signal fork81_outs_0_valid : std_logic;
  signal fork81_outs_0_ready : std_logic;
  signal fork81_outs_1 : std_logic_vector(31 downto 0);
  signal fork81_outs_1_valid : std_logic;
  signal fork81_outs_1_ready : std_logic;
  signal fork81_outs_2 : std_logic_vector(31 downto 0);
  signal fork81_outs_2_valid : std_logic;
  signal fork81_outs_2_ready : std_logic;
  signal mux16_outs : std_logic_vector(4 downto 0);
  signal mux16_outs_valid : std_logic;
  signal mux16_outs_ready : std_logic;
  signal buffer218_outs : std_logic_vector(4 downto 0);
  signal buffer218_outs_valid : std_logic;
  signal buffer218_outs_ready : std_logic;
  signal buffer220_outs : std_logic_vector(4 downto 0);
  signal buffer220_outs_valid : std_logic;
  signal buffer220_outs_ready : std_logic;
  signal fork82_outs_0 : std_logic_vector(4 downto 0);
  signal fork82_outs_0_valid : std_logic;
  signal fork82_outs_0_ready : std_logic;
  signal fork82_outs_1 : std_logic_vector(4 downto 0);
  signal fork82_outs_1_valid : std_logic;
  signal fork82_outs_1_ready : std_logic;
  signal extsi90_outs : std_logic_vector(31 downto 0);
  signal extsi90_outs_valid : std_logic;
  signal extsi90_outs_ready : std_logic;
  signal buffer181_outs : std_logic_vector(4 downto 0);
  signal buffer181_outs_valid : std_logic;
  signal buffer181_outs_ready : std_logic;
  signal fork83_outs_0 : std_logic_vector(31 downto 0);
  signal fork83_outs_0_valid : std_logic;
  signal fork83_outs_0_ready : std_logic;
  signal fork83_outs_1 : std_logic_vector(31 downto 0);
  signal fork83_outs_1_valid : std_logic;
  signal fork83_outs_1_ready : std_logic;
  signal fork83_outs_2 : std_logic_vector(31 downto 0);
  signal fork83_outs_2_valid : std_logic;
  signal fork83_outs_2_ready : std_logic;
  signal fork83_outs_3 : std_logic_vector(31 downto 0);
  signal fork83_outs_3_valid : std_logic;
  signal fork83_outs_3_ready : std_logic;
  signal fork83_outs_4 : std_logic_vector(31 downto 0);
  signal fork83_outs_4_valid : std_logic;
  signal fork83_outs_4_ready : std_logic;
  signal fork83_outs_5 : std_logic_vector(31 downto 0);
  signal fork83_outs_5_valid : std_logic;
  signal fork83_outs_5_ready : std_logic;
  signal mux17_outs : std_logic_vector(4 downto 0);
  signal mux17_outs_valid : std_logic;
  signal mux17_outs_ready : std_logic;
  signal buffer221_outs : std_logic_vector(4 downto 0);
  signal buffer221_outs_valid : std_logic;
  signal buffer221_outs_ready : std_logic;
  signal buffer222_outs : std_logic_vector(4 downto 0);
  signal buffer222_outs_valid : std_logic;
  signal buffer222_outs_ready : std_logic;
  signal fork84_outs_0 : std_logic_vector(4 downto 0);
  signal fork84_outs_0_valid : std_logic;
  signal fork84_outs_0_ready : std_logic;
  signal fork84_outs_1 : std_logic_vector(4 downto 0);
  signal fork84_outs_1_valid : std_logic;
  signal fork84_outs_1_ready : std_logic;
  signal extsi91_outs : std_logic_vector(31 downto 0);
  signal extsi91_outs_valid : std_logic;
  signal extsi91_outs_ready : std_logic;
  signal fork85_outs_0 : std_logic_vector(31 downto 0);
  signal fork85_outs_0_valid : std_logic;
  signal fork85_outs_0_ready : std_logic;
  signal fork85_outs_1 : std_logic_vector(31 downto 0);
  signal fork85_outs_1_valid : std_logic;
  signal fork85_outs_1_ready : std_logic;
  signal fork85_outs_2 : std_logic_vector(31 downto 0);
  signal fork85_outs_2_valid : std_logic;
  signal fork85_outs_2_ready : std_logic;
  signal control_merge12_outs_valid : std_logic;
  signal control_merge12_outs_ready : std_logic;
  signal control_merge12_index : std_logic_vector(0 downto 0);
  signal control_merge12_index_valid : std_logic;
  signal control_merge12_index_ready : std_logic;
  signal fork86_outs_0 : std_logic_vector(0 downto 0);
  signal fork86_outs_0_valid : std_logic;
  signal fork86_outs_0_ready : std_logic;
  signal fork86_outs_1 : std_logic_vector(0 downto 0);
  signal fork86_outs_1_valid : std_logic;
  signal fork86_outs_1_ready : std_logic;
  signal fork86_outs_2 : std_logic_vector(0 downto 0);
  signal fork86_outs_2_valid : std_logic;
  signal fork86_outs_2_ready : std_logic;
  signal buffer224_outs_valid : std_logic;
  signal buffer224_outs_ready : std_logic;
  signal fork87_outs_0_valid : std_logic;
  signal fork87_outs_0_ready : std_logic;
  signal fork87_outs_1_valid : std_logic;
  signal fork87_outs_1_ready : std_logic;
  signal constant79_outs : std_logic_vector(1 downto 0);
  signal constant79_outs_valid : std_logic;
  signal constant79_outs_ready : std_logic;
  signal extsi37_outs : std_logic_vector(31 downto 0);
  signal extsi37_outs_valid : std_logic;
  signal extsi37_outs_ready : std_logic;
  signal source20_outs_valid : std_logic;
  signal source20_outs_ready : std_logic;
  signal constant80_outs : std_logic_vector(4 downto 0);
  signal constant80_outs_valid : std_logic;
  signal constant80_outs_ready : std_logic;
  signal extsi92_outs : std_logic_vector(5 downto 0);
  signal extsi92_outs_valid : std_logic;
  signal extsi92_outs_ready : std_logic;
  signal source21_outs_valid : std_logic;
  signal source21_outs_ready : std_logic;
  signal constant81_outs : std_logic_vector(1 downto 0);
  signal constant81_outs_valid : std_logic;
  signal constant81_outs_ready : std_logic;
  signal fork88_outs_0 : std_logic_vector(1 downto 0);
  signal fork88_outs_0_valid : std_logic;
  signal fork88_outs_0_ready : std_logic;
  signal fork88_outs_1 : std_logic_vector(1 downto 0);
  signal fork88_outs_1_valid : std_logic;
  signal fork88_outs_1_ready : std_logic;
  signal extsi93_outs : std_logic_vector(5 downto 0);
  signal extsi93_outs_valid : std_logic;
  signal extsi93_outs_ready : std_logic;
  signal extsi39_outs : std_logic_vector(31 downto 0);
  signal extsi39_outs_valid : std_logic;
  signal extsi39_outs_ready : std_logic;
  signal buffer185_outs : std_logic_vector(1 downto 0);
  signal buffer185_outs_valid : std_logic;
  signal buffer185_outs_ready : std_logic;
  signal fork89_outs_0 : std_logic_vector(31 downto 0);
  signal fork89_outs_0_valid : std_logic;
  signal fork89_outs_0_ready : std_logic;
  signal fork89_outs_1 : std_logic_vector(31 downto 0);
  signal fork89_outs_1_valid : std_logic;
  signal fork89_outs_1_ready : std_logic;
  signal fork89_outs_2 : std_logic_vector(31 downto 0);
  signal fork89_outs_2_valid : std_logic;
  signal fork89_outs_2_ready : std_logic;
  signal fork89_outs_3 : std_logic_vector(31 downto 0);
  signal fork89_outs_3_valid : std_logic;
  signal fork89_outs_3_ready : std_logic;
  signal source22_outs_valid : std_logic;
  signal source22_outs_ready : std_logic;
  signal constant82_outs : std_logic_vector(2 downto 0);
  signal constant82_outs_valid : std_logic;
  signal constant82_outs_ready : std_logic;
  signal extsi40_outs : std_logic_vector(31 downto 0);
  signal extsi40_outs_valid : std_logic;
  signal extsi40_outs_ready : std_logic;
  signal fork90_outs_0 : std_logic_vector(31 downto 0);
  signal fork90_outs_0_valid : std_logic;
  signal fork90_outs_0_ready : std_logic;
  signal fork90_outs_1 : std_logic_vector(31 downto 0);
  signal fork90_outs_1_valid : std_logic;
  signal fork90_outs_1_ready : std_logic;
  signal fork90_outs_2 : std_logic_vector(31 downto 0);
  signal fork90_outs_2_valid : std_logic;
  signal fork90_outs_2_ready : std_logic;
  signal fork90_outs_3 : std_logic_vector(31 downto 0);
  signal fork90_outs_3_valid : std_logic;
  signal fork90_outs_3_ready : std_logic;
  signal shli22_result : std_logic_vector(31 downto 0);
  signal shli22_result_valid : std_logic;
  signal shli22_result_ready : std_logic;
  signal buffer187_outs : std_logic_vector(31 downto 0);
  signal buffer187_outs_valid : std_logic;
  signal buffer187_outs_ready : std_logic;
  signal shli23_result : std_logic_vector(31 downto 0);
  signal shli23_result_valid : std_logic;
  signal shli23_result_ready : std_logic;
  signal buffer189_outs : std_logic_vector(31 downto 0);
  signal buffer189_outs_valid : std_logic;
  signal buffer189_outs_ready : std_logic;
  signal buffer226_outs : std_logic_vector(31 downto 0);
  signal buffer226_outs_valid : std_logic;
  signal buffer226_outs_ready : std_logic;
  signal buffer227_outs : std_logic_vector(31 downto 0);
  signal buffer227_outs_valid : std_logic;
  signal buffer227_outs_ready : std_logic;
  signal addi38_result : std_logic_vector(31 downto 0);
  signal addi38_result_valid : std_logic;
  signal addi38_result_ready : std_logic;
  signal buffer228_outs : std_logic_vector(31 downto 0);
  signal buffer228_outs_valid : std_logic;
  signal buffer228_outs_ready : std_logic;
  signal addi14_result : std_logic_vector(31 downto 0);
  signal addi14_result_valid : std_logic;
  signal addi14_result_ready : std_logic;
  signal buffer190_outs : std_logic_vector(31 downto 0);
  signal buffer190_outs_valid : std_logic;
  signal buffer190_outs_ready : std_logic;
  signal gate4_outs : std_logic_vector(31 downto 0);
  signal gate4_outs_valid : std_logic;
  signal gate4_outs_ready : std_logic;
  signal trunci24_outs : std_logic_vector(6 downto 0);
  signal trunci24_outs_valid : std_logic;
  signal trunci24_outs_ready : std_logic;
  signal load6_addrOut : std_logic_vector(6 downto 0);
  signal load6_addrOut_valid : std_logic;
  signal load6_addrOut_ready : std_logic;
  signal load6_dataOut : std_logic_vector(31 downto 0);
  signal load6_dataOut_valid : std_logic;
  signal load6_dataOut_ready : std_logic;
  signal shli24_result : std_logic_vector(31 downto 0);
  signal shli24_result_valid : std_logic;
  signal shli24_result_ready : std_logic;
  signal buffer192_outs : std_logic_vector(31 downto 0);
  signal buffer192_outs_valid : std_logic;
  signal buffer192_outs_ready : std_logic;
  signal shli25_result : std_logic_vector(31 downto 0);
  signal shli25_result_valid : std_logic;
  signal shli25_result_ready : std_logic;
  signal buffer194_outs : std_logic_vector(31 downto 0);
  signal buffer194_outs_valid : std_logic;
  signal buffer194_outs_ready : std_logic;
  signal buffer229_outs : std_logic_vector(31 downto 0);
  signal buffer229_outs_valid : std_logic;
  signal buffer229_outs_ready : std_logic;
  signal buffer230_outs : std_logic_vector(31 downto 0);
  signal buffer230_outs_valid : std_logic;
  signal buffer230_outs_ready : std_logic;
  signal addi39_result : std_logic_vector(31 downto 0);
  signal addi39_result_valid : std_logic;
  signal addi39_result_ready : std_logic;
  signal buffer231_outs : std_logic_vector(31 downto 0);
  signal buffer231_outs_valid : std_logic;
  signal buffer231_outs_ready : std_logic;
  signal addi15_result : std_logic_vector(31 downto 0);
  signal addi15_result_valid : std_logic;
  signal addi15_result_ready : std_logic;
  signal gate5_outs : std_logic_vector(31 downto 0);
  signal gate5_outs_valid : std_logic;
  signal gate5_outs_ready : std_logic;
  signal trunci25_outs : std_logic_vector(6 downto 0);
  signal trunci25_outs_valid : std_logic;
  signal trunci25_outs_ready : std_logic;
  signal load7_addrOut : std_logic_vector(6 downto 0);
  signal load7_addrOut_valid : std_logic;
  signal load7_addrOut_ready : std_logic;
  signal load7_dataOut : std_logic_vector(31 downto 0);
  signal load7_dataOut_valid : std_logic;
  signal load7_dataOut_ready : std_logic;
  signal muli2_result : std_logic_vector(31 downto 0);
  signal muli2_result_valid : std_logic;
  signal muli2_result_ready : std_logic;
  signal shli26_result : std_logic_vector(31 downto 0);
  signal shli26_result_valid : std_logic;
  signal shli26_result_ready : std_logic;
  signal buffer196_outs : std_logic_vector(31 downto 0);
  signal buffer196_outs_valid : std_logic;
  signal buffer196_outs_ready : std_logic;
  signal buffer197_outs : std_logic_vector(31 downto 0);
  signal buffer197_outs_valid : std_logic;
  signal buffer197_outs_ready : std_logic;
  signal shli27_result : std_logic_vector(31 downto 0);
  signal shli27_result_valid : std_logic;
  signal shli27_result_ready : std_logic;
  signal buffer198_outs : std_logic_vector(31 downto 0);
  signal buffer198_outs_valid : std_logic;
  signal buffer198_outs_ready : std_logic;
  signal buffer199_outs : std_logic_vector(31 downto 0);
  signal buffer199_outs_valid : std_logic;
  signal buffer199_outs_ready : std_logic;
  signal buffer233_outs : std_logic_vector(31 downto 0);
  signal buffer233_outs_valid : std_logic;
  signal buffer233_outs_ready : std_logic;
  signal buffer234_outs : std_logic_vector(31 downto 0);
  signal buffer234_outs_valid : std_logic;
  signal buffer234_outs_ready : std_logic;
  signal addi40_result : std_logic_vector(31 downto 0);
  signal addi40_result_valid : std_logic;
  signal addi40_result_ready : std_logic;
  signal buffer235_outs : std_logic_vector(31 downto 0);
  signal buffer235_outs_valid : std_logic;
  signal buffer235_outs_ready : std_logic;
  signal addi16_result : std_logic_vector(31 downto 0);
  signal addi16_result_valid : std_logic;
  signal addi16_result_ready : std_logic;
  signal buffer200_outs : std_logic_vector(31 downto 0);
  signal buffer200_outs_valid : std_logic;
  signal buffer200_outs_ready : std_logic;
  signal buffer211_outs_valid : std_logic;
  signal buffer211_outs_ready : std_logic;
  signal gate6_outs : std_logic_vector(31 downto 0);
  signal gate6_outs_valid : std_logic;
  signal gate6_outs_ready : std_logic;
  signal trunci26_outs : std_logic_vector(6 downto 0);
  signal trunci26_outs_valid : std_logic;
  signal trunci26_outs_ready : std_logic;
  signal load8_addrOut : std_logic_vector(6 downto 0);
  signal load8_addrOut_valid : std_logic;
  signal load8_addrOut_ready : std_logic;
  signal load8_dataOut : std_logic_vector(31 downto 0);
  signal load8_dataOut_valid : std_logic;
  signal load8_dataOut_ready : std_logic;
  signal addi2_result : std_logic_vector(31 downto 0);
  signal addi2_result_valid : std_logic;
  signal addi2_result_ready : std_logic;
  signal shli28_result : std_logic_vector(31 downto 0);
  signal shli28_result_valid : std_logic;
  signal shli28_result_ready : std_logic;
  signal buffer201_outs : std_logic_vector(31 downto 0);
  signal buffer201_outs_valid : std_logic;
  signal buffer201_outs_ready : std_logic;
  signal buffer202_outs : std_logic_vector(31 downto 0);
  signal buffer202_outs_valid : std_logic;
  signal buffer202_outs_ready : std_logic;
  signal shli29_result : std_logic_vector(31 downto 0);
  signal shli29_result_valid : std_logic;
  signal shli29_result_ready : std_logic;
  signal buffer203_outs : std_logic_vector(31 downto 0);
  signal buffer203_outs_valid : std_logic;
  signal buffer203_outs_ready : std_logic;
  signal buffer204_outs : std_logic_vector(31 downto 0);
  signal buffer204_outs_valid : std_logic;
  signal buffer204_outs_ready : std_logic;
  signal buffer236_outs : std_logic_vector(31 downto 0);
  signal buffer236_outs_valid : std_logic;
  signal buffer236_outs_ready : std_logic;
  signal buffer237_outs : std_logic_vector(31 downto 0);
  signal buffer237_outs_valid : std_logic;
  signal buffer237_outs_ready : std_logic;
  signal addi41_result : std_logic_vector(31 downto 0);
  signal addi41_result_valid : std_logic;
  signal addi41_result_ready : std_logic;
  signal buffer238_outs : std_logic_vector(31 downto 0);
  signal buffer238_outs_valid : std_logic;
  signal buffer238_outs_ready : std_logic;
  signal addi17_result : std_logic_vector(31 downto 0);
  signal addi17_result_valid : std_logic;
  signal addi17_result_ready : std_logic;
  signal buffer205_outs : std_logic_vector(31 downto 0);
  signal buffer205_outs_valid : std_logic;
  signal buffer205_outs_ready : std_logic;
  signal buffer239_outs_valid : std_logic;
  signal buffer239_outs_ready : std_logic;
  signal buffer5_outs_valid : std_logic;
  signal buffer5_outs_ready : std_logic;
  signal gate7_outs : std_logic_vector(31 downto 0);
  signal gate7_outs_valid : std_logic;
  signal gate7_outs_ready : std_logic;
  signal trunci27_outs : std_logic_vector(6 downto 0);
  signal trunci27_outs_valid : std_logic;
  signal trunci27_outs_ready : std_logic;
  signal store5_addrOut : std_logic_vector(6 downto 0);
  signal store5_addrOut_valid : std_logic;
  signal store5_addrOut_ready : std_logic;
  signal store5_dataToMem : std_logic_vector(31 downto 0);
  signal store5_dataToMem_valid : std_logic;
  signal store5_dataToMem_ready : std_logic;
  signal store5_doneOut_valid : std_logic;
  signal store5_doneOut_ready : std_logic;
  signal addi24_result : std_logic_vector(5 downto 0);
  signal addi24_result_valid : std_logic;
  signal addi24_result_ready : std_logic;
  signal fork91_outs_0 : std_logic_vector(5 downto 0);
  signal fork91_outs_0_valid : std_logic;
  signal fork91_outs_0_ready : std_logic;
  signal fork91_outs_1 : std_logic_vector(5 downto 0);
  signal fork91_outs_1_valid : std_logic;
  signal fork91_outs_1_ready : std_logic;
  signal trunci28_outs : std_logic_vector(4 downto 0);
  signal trunci28_outs_valid : std_logic;
  signal trunci28_outs_ready : std_logic;
  signal buffer206_outs : std_logic_vector(5 downto 0);
  signal buffer206_outs_valid : std_logic;
  signal buffer206_outs_ready : std_logic;
  signal buffer241_outs : std_logic_vector(5 downto 0);
  signal buffer241_outs_valid : std_logic;
  signal buffer241_outs_ready : std_logic;
  signal cmpi6_result : std_logic_vector(0 downto 0);
  signal cmpi6_result_valid : std_logic;
  signal cmpi6_result_ready : std_logic;
  signal buffer207_outs : std_logic_vector(5 downto 0);
  signal buffer207_outs_valid : std_logic;
  signal buffer207_outs_ready : std_logic;
  signal buffer240_outs : std_logic_vector(0 downto 0);
  signal buffer240_outs_valid : std_logic;
  signal buffer240_outs_ready : std_logic;
  signal fork92_outs_0 : std_logic_vector(0 downto 0);
  signal fork92_outs_0_valid : std_logic;
  signal fork92_outs_0_ready : std_logic;
  signal fork92_outs_1 : std_logic_vector(0 downto 0);
  signal fork92_outs_1_valid : std_logic;
  signal fork92_outs_1_ready : std_logic;
  signal fork92_outs_2 : std_logic_vector(0 downto 0);
  signal fork92_outs_2_valid : std_logic;
  signal fork92_outs_2_ready : std_logic;
  signal fork92_outs_3 : std_logic_vector(0 downto 0);
  signal fork92_outs_3_valid : std_logic;
  signal fork92_outs_3_ready : std_logic;
  signal fork92_outs_4 : std_logic_vector(0 downto 0);
  signal fork92_outs_4_valid : std_logic;
  signal fork92_outs_4_ready : std_logic;
  signal fork92_outs_5 : std_logic_vector(0 downto 0);
  signal fork92_outs_5_valid : std_logic;
  signal fork92_outs_5_ready : std_logic;
  signal fork92_outs_6 : std_logic_vector(0 downto 0);
  signal fork92_outs_6_valid : std_logic;
  signal fork92_outs_6_ready : std_logic;
  signal fork92_outs_7 : std_logic_vector(0 downto 0);
  signal fork92_outs_7_valid : std_logic;
  signal fork92_outs_7_ready : std_logic;
  signal fork92_outs_8 : std_logic_vector(0 downto 0);
  signal fork92_outs_8_valid : std_logic;
  signal fork92_outs_8_ready : std_logic;
  signal fork92_outs_9 : std_logic_vector(0 downto 0);
  signal fork92_outs_9_valid : std_logic;
  signal fork92_outs_9_ready : std_logic;
  signal fork92_outs_10 : std_logic_vector(0 downto 0);
  signal fork92_outs_10_valid : std_logic;
  signal fork92_outs_10_ready : std_logic;
  signal cond_br29_trueOut : std_logic_vector(4 downto 0);
  signal cond_br29_trueOut_valid : std_logic;
  signal cond_br29_trueOut_ready : std_logic;
  signal cond_br29_falseOut : std_logic_vector(4 downto 0);
  signal cond_br29_falseOut_valid : std_logic;
  signal cond_br29_falseOut_ready : std_logic;
  signal cond_br30_trueOut : std_logic_vector(4 downto 0);
  signal cond_br30_trueOut_valid : std_logic;
  signal cond_br30_trueOut_ready : std_logic;
  signal cond_br30_falseOut : std_logic_vector(4 downto 0);
  signal cond_br30_falseOut_valid : std_logic;
  signal cond_br30_falseOut_ready : std_logic;
  signal buffer209_outs : std_logic_vector(0 downto 0);
  signal buffer209_outs_valid : std_logic;
  signal buffer209_outs_ready : std_logic;
  signal buffer210_outs : std_logic_vector(4 downto 0);
  signal buffer210_outs_valid : std_logic;
  signal buffer210_outs_ready : std_logic;
  signal cond_br31_trueOut : std_logic_vector(4 downto 0);
  signal cond_br31_trueOut_valid : std_logic;
  signal cond_br31_trueOut_ready : std_logic;
  signal cond_br31_falseOut : std_logic_vector(4 downto 0);
  signal cond_br31_falseOut_valid : std_logic;
  signal cond_br31_falseOut_ready : std_logic;
  signal buffer212_outs : std_logic_vector(4 downto 0);
  signal buffer212_outs_valid : std_logic;
  signal buffer212_outs_ready : std_logic;
  signal cond_br32_trueOut_valid : std_logic;
  signal cond_br32_trueOut_ready : std_logic;
  signal cond_br32_falseOut_valid : std_logic;
  signal cond_br32_falseOut_ready : std_logic;
  signal buffer213_outs : std_logic_vector(0 downto 0);
  signal buffer213_outs_valid : std_logic;
  signal buffer213_outs_ready : std_logic;
  signal cond_br134_trueOut_valid : std_logic;
  signal cond_br134_trueOut_ready : std_logic;
  signal cond_br134_falseOut_valid : std_logic;
  signal cond_br134_falseOut_ready : std_logic;
  signal buffer214_outs : std_logic_vector(0 downto 0);
  signal buffer214_outs_valid : std_logic;
  signal buffer214_outs_ready : std_logic;
  signal cond_br135_trueOut_valid : std_logic;
  signal cond_br135_trueOut_ready : std_logic;
  signal cond_br135_falseOut_valid : std_logic;
  signal cond_br135_falseOut_ready : std_logic;
  signal cond_br136_trueOut_valid : std_logic;
  signal cond_br136_trueOut_ready : std_logic;
  signal cond_br136_falseOut_valid : std_logic;
  signal cond_br136_falseOut_ready : std_logic;
  signal cond_br137_trueOut_valid : std_logic;
  signal cond_br137_trueOut_ready : std_logic;
  signal cond_br137_falseOut_valid : std_logic;
  signal cond_br137_falseOut_ready : std_logic;
  signal buffer217_outs : std_logic_vector(0 downto 0);
  signal buffer217_outs_valid : std_logic;
  signal buffer217_outs_ready : std_logic;
  signal cond_br138_trueOut_valid : std_logic;
  signal cond_br138_trueOut_ready : std_logic;
  signal cond_br138_falseOut_valid : std_logic;
  signal cond_br138_falseOut_ready : std_logic;
  signal extsi94_outs : std_logic_vector(5 downto 0);
  signal extsi94_outs_valid : std_logic;
  signal extsi94_outs_ready : std_logic;
  signal source23_outs_valid : std_logic;
  signal source23_outs_ready : std_logic;
  signal constant83_outs : std_logic_vector(4 downto 0);
  signal constant83_outs_valid : std_logic;
  signal constant83_outs_ready : std_logic;
  signal extsi95_outs : std_logic_vector(5 downto 0);
  signal extsi95_outs_valid : std_logic;
  signal extsi95_outs_ready : std_logic;
  signal source24_outs_valid : std_logic;
  signal source24_outs_ready : std_logic;
  signal constant84_outs : std_logic_vector(1 downto 0);
  signal constant84_outs_valid : std_logic;
  signal constant84_outs_ready : std_logic;
  signal extsi96_outs : std_logic_vector(5 downto 0);
  signal extsi96_outs_valid : std_logic;
  signal extsi96_outs_ready : std_logic;
  signal addi25_result : std_logic_vector(5 downto 0);
  signal addi25_result_valid : std_logic;
  signal addi25_result_ready : std_logic;
  signal buffer243_outs : std_logic_vector(5 downto 0);
  signal buffer243_outs_valid : std_logic;
  signal buffer243_outs_ready : std_logic;
  signal fork93_outs_0 : std_logic_vector(5 downto 0);
  signal fork93_outs_0_valid : std_logic;
  signal fork93_outs_0_ready : std_logic;
  signal fork93_outs_1 : std_logic_vector(5 downto 0);
  signal fork93_outs_1_valid : std_logic;
  signal fork93_outs_1_ready : std_logic;
  signal trunci29_outs : std_logic_vector(4 downto 0);
  signal trunci29_outs_valid : std_logic;
  signal trunci29_outs_ready : std_logic;
  signal buffer219_outs : std_logic_vector(5 downto 0);
  signal buffer219_outs_valid : std_logic;
  signal buffer219_outs_ready : std_logic;
  signal cmpi7_result : std_logic_vector(0 downto 0);
  signal cmpi7_result_valid : std_logic;
  signal cmpi7_result_ready : std_logic;
  signal buffer244_outs : std_logic_vector(0 downto 0);
  signal buffer244_outs_valid : std_logic;
  signal buffer244_outs_ready : std_logic;
  signal fork94_outs_0 : std_logic_vector(0 downto 0);
  signal fork94_outs_0_valid : std_logic;
  signal fork94_outs_0_ready : std_logic;
  signal fork94_outs_1 : std_logic_vector(0 downto 0);
  signal fork94_outs_1_valid : std_logic;
  signal fork94_outs_1_ready : std_logic;
  signal fork94_outs_2 : std_logic_vector(0 downto 0);
  signal fork94_outs_2_valid : std_logic;
  signal fork94_outs_2_ready : std_logic;
  signal fork94_outs_3 : std_logic_vector(0 downto 0);
  signal fork94_outs_3_valid : std_logic;
  signal fork94_outs_3_ready : std_logic;
  signal fork94_outs_4 : std_logic_vector(0 downto 0);
  signal fork94_outs_4_valid : std_logic;
  signal fork94_outs_4_ready : std_logic;
  signal fork94_outs_5 : std_logic_vector(0 downto 0);
  signal fork94_outs_5_valid : std_logic;
  signal fork94_outs_5_ready : std_logic;
  signal fork94_outs_6 : std_logic_vector(0 downto 0);
  signal fork94_outs_6_valid : std_logic;
  signal fork94_outs_6_ready : std_logic;
  signal fork94_outs_7 : std_logic_vector(0 downto 0);
  signal fork94_outs_7_valid : std_logic;
  signal fork94_outs_7_ready : std_logic;
  signal fork94_outs_8 : std_logic_vector(0 downto 0);
  signal fork94_outs_8_valid : std_logic;
  signal fork94_outs_8_ready : std_logic;
  signal cond_br33_trueOut : std_logic_vector(4 downto 0);
  signal cond_br33_trueOut_valid : std_logic;
  signal cond_br33_trueOut_ready : std_logic;
  signal cond_br33_falseOut : std_logic_vector(4 downto 0);
  signal cond_br33_falseOut_valid : std_logic;
  signal cond_br33_falseOut_ready : std_logic;
  signal cond_br34_trueOut : std_logic_vector(4 downto 0);
  signal cond_br34_trueOut_valid : std_logic;
  signal cond_br34_trueOut_ready : std_logic;
  signal cond_br34_falseOut : std_logic_vector(4 downto 0);
  signal cond_br34_falseOut_valid : std_logic;
  signal cond_br34_falseOut_ready : std_logic;
  signal cond_br35_trueOut_valid : std_logic;
  signal cond_br35_trueOut_ready : std_logic;
  signal cond_br35_falseOut_valid : std_logic;
  signal cond_br35_falseOut_ready : std_logic;
  signal buffer223_outs : std_logic_vector(0 downto 0);
  signal buffer223_outs_valid : std_logic;
  signal buffer223_outs_ready : std_logic;
  signal cond_br139_trueOut_valid : std_logic;
  signal cond_br139_trueOut_ready : std_logic;
  signal cond_br139_falseOut_valid : std_logic;
  signal cond_br139_falseOut_ready : std_logic;
  signal cond_br140_trueOut_valid : std_logic;
  signal cond_br140_trueOut_ready : std_logic;
  signal cond_br140_falseOut_valid : std_logic;
  signal cond_br140_falseOut_ready : std_logic;
  signal buffer225_outs : std_logic_vector(0 downto 0);
  signal buffer225_outs_valid : std_logic;
  signal buffer225_outs_ready : std_logic;
  signal cond_br141_trueOut_valid : std_logic;
  signal cond_br141_trueOut_ready : std_logic;
  signal cond_br141_falseOut_valid : std_logic;
  signal cond_br141_falseOut_ready : std_logic;
  signal cond_br142_trueOut_valid : std_logic;
  signal cond_br142_trueOut_ready : std_logic;
  signal cond_br142_falseOut_valid : std_logic;
  signal cond_br142_falseOut_ready : std_logic;
  signal cond_br143_trueOut_valid : std_logic;
  signal cond_br143_trueOut_ready : std_logic;
  signal cond_br143_falseOut_valid : std_logic;
  signal cond_br143_falseOut_ready : std_logic;
  signal buffer246_outs : std_logic_vector(4 downto 0);
  signal buffer246_outs_valid : std_logic;
  signal buffer246_outs_ready : std_logic;
  signal extsi97_outs : std_logic_vector(5 downto 0);
  signal extsi97_outs_valid : std_logic;
  signal extsi97_outs_ready : std_logic;
  signal source25_outs_valid : std_logic;
  signal source25_outs_ready : std_logic;
  signal constant85_outs : std_logic_vector(4 downto 0);
  signal constant85_outs_valid : std_logic;
  signal constant85_outs_ready : std_logic;
  signal extsi98_outs : std_logic_vector(5 downto 0);
  signal extsi98_outs_valid : std_logic;
  signal extsi98_outs_ready : std_logic;
  signal source26_outs_valid : std_logic;
  signal source26_outs_ready : std_logic;
  signal constant86_outs : std_logic_vector(1 downto 0);
  signal constant86_outs_valid : std_logic;
  signal constant86_outs_ready : std_logic;
  signal extsi99_outs : std_logic_vector(5 downto 0);
  signal extsi99_outs_valid : std_logic;
  signal extsi99_outs_ready : std_logic;
  signal addi26_result : std_logic_vector(5 downto 0);
  signal addi26_result_valid : std_logic;
  signal addi26_result_ready : std_logic;
  signal buffer247_outs : std_logic_vector(5 downto 0);
  signal buffer247_outs_valid : std_logic;
  signal buffer247_outs_ready : std_logic;
  signal fork95_outs_0 : std_logic_vector(5 downto 0);
  signal fork95_outs_0_valid : std_logic;
  signal fork95_outs_0_ready : std_logic;
  signal fork95_outs_1 : std_logic_vector(5 downto 0);
  signal fork95_outs_1_valid : std_logic;
  signal fork95_outs_1_ready : std_logic;
  signal trunci30_outs : std_logic_vector(4 downto 0);
  signal trunci30_outs_valid : std_logic;
  signal trunci30_outs_ready : std_logic;
  signal cmpi8_result : std_logic_vector(0 downto 0);
  signal cmpi8_result_valid : std_logic;
  signal cmpi8_result_ready : std_logic;
  signal buffer248_outs : std_logic_vector(0 downto 0);
  signal buffer248_outs_valid : std_logic;
  signal buffer248_outs_ready : std_logic;
  signal fork96_outs_0 : std_logic_vector(0 downto 0);
  signal fork96_outs_0_valid : std_logic;
  signal fork96_outs_0_ready : std_logic;
  signal fork96_outs_1 : std_logic_vector(0 downto 0);
  signal fork96_outs_1_valid : std_logic;
  signal fork96_outs_1_ready : std_logic;
  signal fork96_outs_2 : std_logic_vector(0 downto 0);
  signal fork96_outs_2_valid : std_logic;
  signal fork96_outs_2_ready : std_logic;
  signal fork96_outs_3 : std_logic_vector(0 downto 0);
  signal fork96_outs_3_valid : std_logic;
  signal fork96_outs_3_ready : std_logic;
  signal fork96_outs_4 : std_logic_vector(0 downto 0);
  signal fork96_outs_4_valid : std_logic;
  signal fork96_outs_4_ready : std_logic;
  signal fork96_outs_5 : std_logic_vector(0 downto 0);
  signal fork96_outs_5_valid : std_logic;
  signal fork96_outs_5_ready : std_logic;
  signal fork96_outs_6 : std_logic_vector(0 downto 0);
  signal fork96_outs_6_valid : std_logic;
  signal fork96_outs_6_ready : std_logic;
  signal fork96_outs_7 : std_logic_vector(0 downto 0);
  signal fork96_outs_7_valid : std_logic;
  signal fork96_outs_7_ready : std_logic;
  signal cond_br36_trueOut : std_logic_vector(4 downto 0);
  signal cond_br36_trueOut_valid : std_logic;
  signal cond_br36_trueOut_ready : std_logic;
  signal cond_br36_falseOut : std_logic_vector(4 downto 0);
  signal cond_br36_falseOut_valid : std_logic;
  signal cond_br36_falseOut_ready : std_logic;
  signal cond_br37_trueOut_valid : std_logic;
  signal cond_br37_trueOut_ready : std_logic;
  signal cond_br37_falseOut_valid : std_logic;
  signal cond_br37_falseOut_ready : std_logic;
  signal buffer232_outs : std_logic_vector(0 downto 0);
  signal buffer232_outs_valid : std_logic;
  signal buffer232_outs_ready : std_logic;
  signal fork97_outs_0_valid : std_logic;
  signal fork97_outs_0_ready : std_logic;
  signal fork97_outs_1_valid : std_logic;
  signal fork97_outs_1_ready : std_logic;
  signal fork97_outs_2_valid : std_logic;
  signal fork97_outs_2_ready : std_logic;
  signal fork97_outs_3_valid : std_logic;
  signal fork97_outs_3_ready : std_logic;
  signal fork97_outs_4_valid : std_logic;
  signal fork97_outs_4_ready : std_logic;
  signal fork97_outs_5_valid : std_logic;
  signal fork97_outs_5_ready : std_logic;
  signal fork97_outs_6_valid : std_logic;
  signal fork97_outs_6_ready : std_logic;

begin

  A_end_valid <= mem_controller10_memEnd_valid;
  mem_controller10_memEnd_ready <= A_end_ready;
  B_end_valid <= mem_controller9_memEnd_valid;
  mem_controller9_memEnd_ready <= B_end_ready;
  C_end_valid <= mem_controller8_memEnd_valid;
  mem_controller8_memEnd_ready <= C_end_ready;
  D_end_valid <= mem_controller7_memEnd_valid;
  mem_controller7_memEnd_ready <= D_end_ready;
  E_end_valid <= mem_controller6_memEnd_valid;
  mem_controller6_memEnd_ready <= E_end_ready;
  F_end_valid <= mem_controller5_memEnd_valid;
  mem_controller5_memEnd_ready <= F_end_ready;
  G_end_valid <= mem_controller4_memEnd_valid;
  mem_controller4_memEnd_ready <= G_end_ready;
  end_valid <= fork0_outs_1_valid;
  fork0_outs_1_ready <= end_ready;
  A_loadEn <= mem_controller10_loadEn;
  A_loadAddr <= mem_controller10_loadAddr;
  A_storeEn <= mem_controller10_storeEn;
  A_storeAddr <= mem_controller10_storeAddr;
  A_storeData <= mem_controller10_storeData;
  B_loadEn <= mem_controller9_loadEn;
  B_loadAddr <= mem_controller9_loadAddr;
  B_storeEn <= mem_controller9_storeEn;
  B_storeAddr <= mem_controller9_storeAddr;
  B_storeData <= mem_controller9_storeData;
  C_loadEn <= mem_controller8_loadEn;
  C_loadAddr <= mem_controller8_loadAddr;
  C_storeEn <= mem_controller8_storeEn;
  C_storeAddr <= mem_controller8_storeAddr;
  C_storeData <= mem_controller8_storeData;
  D_loadEn <= mem_controller7_loadEn;
  D_loadAddr <= mem_controller7_loadAddr;
  D_storeEn <= mem_controller7_storeEn;
  D_storeAddr <= mem_controller7_storeAddr;
  D_storeData <= mem_controller7_storeData;
  E_loadEn <= mem_controller6_loadEn;
  E_loadAddr <= mem_controller6_loadAddr;
  E_storeEn <= mem_controller6_storeEn;
  E_storeAddr <= mem_controller6_storeAddr;
  E_storeData <= mem_controller6_storeData;
  F_loadEn <= mem_controller5_loadEn;
  F_loadAddr <= mem_controller5_loadAddr;
  F_storeEn <= mem_controller5_storeEn;
  F_storeAddr <= mem_controller5_storeAddr;
  F_storeData <= mem_controller5_storeData;
  G_loadEn <= mem_controller4_loadEn;
  G_loadAddr <= mem_controller4_loadAddr;
  G_storeEn <= mem_controller4_storeEn;
  G_storeAddr <= mem_controller4_storeAddr;
  G_storeData <= mem_controller4_storeData;

  fork0 : entity work.fork_dataless(arch) generic map(6)
    port map(
      ins_valid => start_valid,
      ins_ready => start_ready,
      clk => clk,
      rst => rst,
      outs_valid(0) => fork0_outs_0_valid,
      outs_valid(1) => fork0_outs_1_valid,
      outs_valid(2) => fork0_outs_2_valid,
      outs_valid(3) => fork0_outs_3_valid,
      outs_valid(4) => fork0_outs_4_valid,
      outs_valid(5) => fork0_outs_5_valid,
      outs_ready(0) => fork0_outs_0_ready,
      outs_ready(1) => fork0_outs_1_ready,
      outs_ready(2) => fork0_outs_2_ready,
      outs_ready(3) => fork0_outs_3_ready,
      outs_ready(4) => fork0_outs_4_ready,
      outs_ready(5) => fork0_outs_5_ready
    );

  mem_controller4 : entity work.mem_controller(arch) generic map(2, 1, 2, 32, 7)
    port map(
      loadData => G_loadData,
      memStart_valid => G_start_valid,
      memStart_ready => G_start_ready,
      ctrl(0) => extsi32_outs,
      ctrl(1) => extsi37_outs,
      ctrl_valid(0) => extsi32_outs_valid,
      ctrl_valid(1) => extsi37_outs_valid,
      ctrl_ready(0) => extsi32_outs_ready,
      ctrl_ready(1) => extsi37_outs_ready,
      stAddr(0) => store4_addrOut,
      stAddr(1) => store5_addrOut,
      stAddr_valid(0) => store4_addrOut_valid,
      stAddr_valid(1) => store5_addrOut_valid,
      stAddr_ready(0) => store4_addrOut_ready,
      stAddr_ready(1) => store5_addrOut_ready,
      stData(0) => store4_dataToMem,
      stData(1) => store5_dataToMem,
      stData_valid(0) => store4_dataToMem_valid,
      stData_valid(1) => store5_dataToMem_valid,
      stData_ready(0) => store4_dataToMem_ready,
      stData_ready(1) => store5_dataToMem_ready,
      ldAddr(0) => load8_addrOut,
      ldAddr_valid(0) => load8_addrOut_valid,
      ldAddr_ready(0) => load8_addrOut_ready,
      ctrlEnd_valid => fork97_outs_6_valid,
      ctrlEnd_ready => fork97_outs_6_ready,
      clk => clk,
      rst => rst,
      stDone_valid(0) => mem_controller4_stDone_0_valid,
      stDone_valid(1) => mem_controller4_stDone_1_valid,
      stDone_ready(0) => mem_controller4_stDone_0_ready,
      stDone_ready(1) => mem_controller4_stDone_1_ready,
      ldData(0) => mem_controller4_ldData_0,
      ldData_valid(0) => mem_controller4_ldData_0_valid,
      ldData_ready(0) => mem_controller4_ldData_0_ready,
      memEnd_valid => mem_controller4_memEnd_valid,
      memEnd_ready => mem_controller4_memEnd_ready,
      loadEn => mem_controller4_loadEn,
      loadAddr => mem_controller4_loadAddr,
      storeEn => mem_controller4_storeEn,
      storeAddr => mem_controller4_storeAddr,
      storeData => mem_controller4_storeData
    );

  mem_controller5 : entity work.mem_controller(arch) generic map(2, 2, 2, 32, 7)
    port map(
      loadData => F_loadData,
      memStart_valid => F_start_valid,
      memStart_ready => F_start_ready,
      ctrl(0) => extsi17_outs,
      ctrl(1) => extsi22_outs,
      ctrl_valid(0) => extsi17_outs_valid,
      ctrl_valid(1) => extsi22_outs_valid,
      ctrl_ready(0) => extsi17_outs_ready,
      ctrl_ready(1) => extsi22_outs_ready,
      stAddr(0) => store2_addrOut,
      stAddr(1) => store3_addrOut,
      stAddr_valid(0) => store2_addrOut_valid,
      stAddr_valid(1) => store3_addrOut_valid,
      stAddr_ready(0) => store2_addrOut_ready,
      stAddr_ready(1) => store3_addrOut_ready,
      stData(0) => store2_dataToMem,
      stData(1) => store3_dataToMem,
      stData_valid(0) => store2_dataToMem_valid,
      stData_valid(1) => store3_dataToMem_valid,
      stData_ready(0) => store2_dataToMem_ready,
      stData_ready(1) => store3_dataToMem_ready,
      ldAddr(0) => load5_addrOut,
      ldAddr(1) => load7_addrOut,
      ldAddr_valid(0) => load5_addrOut_valid,
      ldAddr_valid(1) => load7_addrOut_valid,
      ldAddr_ready(0) => load5_addrOut_ready,
      ldAddr_ready(1) => load7_addrOut_ready,
      ctrlEnd_valid => fork97_outs_5_valid,
      ctrlEnd_ready => fork97_outs_5_ready,
      clk => clk,
      rst => rst,
      stDone_valid(0) => mem_controller5_stDone_0_valid,
      stDone_valid(1) => mem_controller5_stDone_1_valid,
      stDone_ready(0) => mem_controller5_stDone_0_ready,
      stDone_ready(1) => mem_controller5_stDone_1_ready,
      ldData(0) => mem_controller5_ldData_0,
      ldData(1) => mem_controller5_ldData_1,
      ldData_valid(0) => mem_controller5_ldData_0_valid,
      ldData_valid(1) => mem_controller5_ldData_1_valid,
      ldData_ready(0) => mem_controller5_ldData_0_ready,
      ldData_ready(1) => mem_controller5_ldData_1_ready,
      memEnd_valid => mem_controller5_memEnd_valid,
      memEnd_ready => mem_controller5_memEnd_ready,
      loadEn => mem_controller5_loadEn,
      loadAddr => mem_controller5_loadAddr,
      storeEn => mem_controller5_storeEn,
      storeAddr => mem_controller5_storeAddr,
      storeData => mem_controller5_storeData
    );

  mem_controller6 : entity work.mem_controller(arch) generic map(2, 2, 2, 32, 7)
    port map(
      loadData => E_loadData,
      memStart_valid => E_start_valid,
      memStart_ready => E_start_ready,
      ctrl(0) => extsi2_outs,
      ctrl(1) => extsi7_outs,
      ctrl_valid(0) => extsi2_outs_valid,
      ctrl_valid(1) => extsi7_outs_valid,
      ctrl_ready(0) => extsi2_outs_ready,
      ctrl_ready(1) => extsi7_outs_ready,
      stAddr(0) => store0_addrOut,
      stAddr(1) => store1_addrOut,
      stAddr_valid(0) => store0_addrOut_valid,
      stAddr_valid(1) => store1_addrOut_valid,
      stAddr_ready(0) => store0_addrOut_ready,
      stAddr_ready(1) => store1_addrOut_ready,
      stData(0) => store0_dataToMem,
      stData(1) => store1_dataToMem,
      stData_valid(0) => store0_dataToMem_valid,
      stData_valid(1) => store1_dataToMem_valid,
      stData_ready(0) => store0_dataToMem_ready,
      stData_ready(1) => store1_dataToMem_ready,
      ldAddr(0) => load2_addrOut,
      ldAddr(1) => load6_addrOut,
      ldAddr_valid(0) => load2_addrOut_valid,
      ldAddr_valid(1) => load6_addrOut_valid,
      ldAddr_ready(0) => load2_addrOut_ready,
      ldAddr_ready(1) => load6_addrOut_ready,
      ctrlEnd_valid => fork97_outs_4_valid,
      ctrlEnd_ready => fork97_outs_4_ready,
      clk => clk,
      rst => rst,
      stDone_valid(0) => mem_controller6_stDone_0_valid,
      stDone_valid(1) => mem_controller6_stDone_1_valid,
      stDone_ready(0) => mem_controller6_stDone_0_ready,
      stDone_ready(1) => mem_controller6_stDone_1_ready,
      ldData(0) => mem_controller6_ldData_0,
      ldData(1) => mem_controller6_ldData_1,
      ldData_valid(0) => mem_controller6_ldData_0_valid,
      ldData_valid(1) => mem_controller6_ldData_1_valid,
      ldData_ready(0) => mem_controller6_ldData_0_ready,
      ldData_ready(1) => mem_controller6_ldData_1_ready,
      memEnd_valid => mem_controller6_memEnd_valid,
      memEnd_ready => mem_controller6_memEnd_ready,
      loadEn => mem_controller6_loadEn,
      loadAddr => mem_controller6_loadAddr,
      storeEn => mem_controller6_storeEn,
      storeAddr => mem_controller6_storeAddr,
      storeData => mem_controller6_storeData
    );

  mem_controller7 : entity work.mem_controller_storeless(arch) generic map(1, 32, 7)
    port map(
      loadData => D_loadData,
      memStart_valid => D_start_valid,
      memStart_ready => D_start_ready,
      ldAddr(0) => load4_addrOut,
      ldAddr_valid(0) => load4_addrOut_valid,
      ldAddr_ready(0) => load4_addrOut_ready,
      ctrlEnd_valid => fork97_outs_3_valid,
      ctrlEnd_ready => fork97_outs_3_ready,
      clk => clk,
      rst => rst,
      ldData(0) => mem_controller7_ldData_0,
      ldData_valid(0) => mem_controller7_ldData_0_valid,
      ldData_ready(0) => mem_controller7_ldData_0_ready,
      memEnd_valid => mem_controller7_memEnd_valid,
      memEnd_ready => mem_controller7_memEnd_ready,
      loadEn => mem_controller7_loadEn,
      loadAddr => mem_controller7_loadAddr,
      storeEn => mem_controller7_storeEn,
      storeAddr => mem_controller7_storeAddr,
      storeData => mem_controller7_storeData
    );

  mem_controller8 : entity work.mem_controller_storeless(arch) generic map(1, 32, 7)
    port map(
      loadData => C_loadData,
      memStart_valid => C_start_valid,
      memStart_ready => C_start_ready,
      ldAddr(0) => load3_addrOut,
      ldAddr_valid(0) => load3_addrOut_valid,
      ldAddr_ready(0) => load3_addrOut_ready,
      ctrlEnd_valid => fork97_outs_2_valid,
      ctrlEnd_ready => fork97_outs_2_ready,
      clk => clk,
      rst => rst,
      ldData(0) => mem_controller8_ldData_0,
      ldData_valid(0) => mem_controller8_ldData_0_valid,
      ldData_ready(0) => mem_controller8_ldData_0_ready,
      memEnd_valid => mem_controller8_memEnd_valid,
      memEnd_ready => mem_controller8_memEnd_ready,
      loadEn => mem_controller8_loadEn,
      loadAddr => mem_controller8_loadAddr,
      storeEn => mem_controller8_storeEn,
      storeAddr => mem_controller8_storeAddr,
      storeData => mem_controller8_storeData
    );

  mem_controller9 : entity work.mem_controller_storeless(arch) generic map(1, 32, 7)
    port map(
      loadData => B_loadData,
      memStart_valid => B_start_valid,
      memStart_ready => B_start_ready,
      ldAddr(0) => load1_addrOut,
      ldAddr_valid(0) => load1_addrOut_valid,
      ldAddr_ready(0) => load1_addrOut_ready,
      ctrlEnd_valid => fork97_outs_1_valid,
      ctrlEnd_ready => fork97_outs_1_ready,
      clk => clk,
      rst => rst,
      ldData(0) => mem_controller9_ldData_0,
      ldData_valid(0) => mem_controller9_ldData_0_valid,
      ldData_ready(0) => mem_controller9_ldData_0_ready,
      memEnd_valid => mem_controller9_memEnd_valid,
      memEnd_ready => mem_controller9_memEnd_ready,
      loadEn => mem_controller9_loadEn,
      loadAddr => mem_controller9_loadAddr,
      storeEn => mem_controller9_storeEn,
      storeAddr => mem_controller9_storeAddr,
      storeData => mem_controller9_storeData
    );

  mem_controller10 : entity work.mem_controller_storeless(arch) generic map(1, 32, 7)
    port map(
      loadData => A_loadData,
      memStart_valid => A_start_valid,
      memStart_ready => A_start_ready,
      ldAddr(0) => load0_addrOut,
      ldAddr_valid(0) => load0_addrOut_valid,
      ldAddr_ready(0) => load0_addrOut_ready,
      ctrlEnd_valid => fork97_outs_0_valid,
      ctrlEnd_ready => fork97_outs_0_ready,
      clk => clk,
      rst => rst,
      ldData(0) => mem_controller10_ldData_0,
      ldData_valid(0) => mem_controller10_ldData_0_valid,
      ldData_ready(0) => mem_controller10_ldData_0_ready,
      memEnd_valid => mem_controller10_memEnd_valid,
      memEnd_ready => mem_controller10_memEnd_ready,
      loadEn => mem_controller10_loadEn,
      loadAddr => mem_controller10_loadAddr,
      storeEn => mem_controller10_storeEn,
      storeAddr => mem_controller10_storeAddr,
      storeData => mem_controller10_storeData
    );

  constant45 : entity work.handshake_constant_0(arch) generic map(1)
    port map(
      ctrl_valid => fork0_outs_0_valid,
      ctrl_ready => fork0_outs_0_ready,
      clk => clk,
      rst => rst,
      outs => constant45_outs,
      outs_valid => constant45_outs_valid,
      outs_ready => constant45_outs_ready
    );

  extsi53 : entity work.extsi(arch) generic map(1, 5)
    port map(
      ins => constant45_outs,
      ins_valid => constant45_outs_valid,
      ins_ready => constant45_outs_ready,
      clk => clk,
      rst => rst,
      outs => extsi53_outs,
      outs_valid => extsi53_outs_valid,
      outs_ready => extsi53_outs_ready
    );

  mux22 : entity work.mux_dataless(arch) generic map(2, 1)
    port map(
      index => init0_outs,
      index_valid => init0_outs_valid,
      index_ready => init0_outs_ready,
      ins_valid(0) => fork0_outs_4_valid,
      ins_valid(1) => cond_br120_trueOut_valid,
      ins_ready(0) => fork0_outs_4_ready,
      ins_ready(1) => cond_br120_trueOut_ready,
      clk => clk,
      rst => rst,
      outs_valid => mux22_outs_valid,
      outs_ready => mux22_outs_ready
    );

  init0 : entity work.tehb_init(arch) generic map(1, 0)
    port map(
      ins => fork28_outs_3,
      ins_valid => fork28_outs_3_valid,
      ins_ready => fork28_outs_3_ready,
      clk => clk,
      rst => rst,
      outs => init0_outs,
      outs_valid => init0_outs_valid,
      outs_ready => init0_outs_ready
    );

  mux0 : entity work.mux(arch) generic map(2, 5, 1)
    port map(
      index => control_merge0_index,
      index_valid => control_merge0_index_valid,
      index_ready => control_merge0_index_ready,
      ins(0) => extsi53_outs,
      ins(1) => cond_br16_trueOut,
      ins_valid(0) => extsi53_outs_valid,
      ins_valid(1) => cond_br16_trueOut_valid,
      ins_ready(0) => extsi53_outs_ready,
      ins_ready(1) => cond_br16_trueOut_ready,
      clk => clk,
      rst => rst,
      outs => mux0_outs,
      outs_valid => mux0_outs_valid,
      outs_ready => mux0_outs_ready
    );

  control_merge0 : entity work.control_merge_dataless(arch) generic map(2, 1)
    port map(
      ins_valid(0) => fork0_outs_5_valid,
      ins_valid(1) => cond_br17_trueOut_valid,
      ins_ready(0) => fork0_outs_5_ready,
      ins_ready(1) => cond_br17_trueOut_ready,
      clk => clk,
      rst => rst,
      outs_valid => control_merge0_outs_valid,
      outs_ready => control_merge0_outs_ready,
      index => control_merge0_index,
      index_valid => control_merge0_index_valid,
      index_ready => control_merge0_index_ready
    );

  fork1 : entity work.fork_dataless(arch) generic map(2)
    port map(
      ins_valid => control_merge0_outs_valid,
      ins_ready => control_merge0_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid(0) => fork1_outs_0_valid,
      outs_valid(1) => fork1_outs_1_valid,
      outs_ready(0) => fork1_outs_0_ready,
      outs_ready(1) => fork1_outs_1_ready
    );

  constant46 : entity work.handshake_constant_0(arch) generic map(1)
    port map(
      ctrl_valid => fork1_outs_0_valid,
      ctrl_ready => fork1_outs_0_ready,
      clk => clk,
      rst => rst,
      outs => constant46_outs,
      outs_valid => constant46_outs_valid,
      outs_ready => constant46_outs_ready
    );

  extsi52 : entity work.extsi(arch) generic map(1, 5)
    port map(
      ins => constant46_outs,
      ins_valid => constant46_outs_valid,
      ins_ready => constant46_outs_ready,
      clk => clk,
      rst => rst,
      outs => extsi52_outs,
      outs_valid => extsi52_outs_valid,
      outs_ready => extsi52_outs_ready
    );

  buffer8 : entity work.tehb(arch) generic map(5)
    port map(
      ins => mux0_outs,
      ins_valid => mux0_outs_valid,
      ins_ready => mux0_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer8_outs,
      outs_valid => buffer8_outs_valid,
      outs_ready => buffer8_outs_ready
    );

  buffer6 : entity work.tehb_dataless(arch)
    port map(
      ins_valid => mux22_outs_valid,
      ins_ready => mux22_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer6_outs_valid,
      outs_ready => buffer6_outs_ready
    );

  mux27 : entity work.mux_dataless(arch) generic map(2, 1)
    port map(
      index => init5_outs,
      index_valid => init5_outs_valid,
      index_ready => init5_outs_ready,
      ins_valid(0) => buffer6_outs_valid,
      ins_valid(1) => cond_br118_trueOut_valid,
      ins_ready(0) => buffer6_outs_ready,
      ins_ready(1) => cond_br118_trueOut_ready,
      clk => clk,
      rst => rst,
      outs_valid => mux27_outs_valid,
      outs_ready => mux27_outs_ready
    );

  init5 : entity work.tehb_init(arch) generic map(1, 0)
    port map(
      ins => buffer7_outs,
      ins_valid => buffer7_outs_valid,
      ins_ready => buffer7_outs_ready,
      clk => clk,
      rst => rst,
      outs => init5_outs,
      outs_valid => init5_outs_valid,
      outs_ready => init5_outs_ready
    );

  buffer7 : entity work.tfifo(arch) generic map(1, 1)
    port map(
      ins => fork25_outs_4,
      ins_valid => fork25_outs_4_valid,
      ins_ready => fork25_outs_4_ready,
      clk => clk,
      rst => rst,
      outs => buffer7_outs,
      outs_valid => buffer7_outs_valid,
      outs_ready => buffer7_outs_ready
    );

  mux1 : entity work.mux(arch) generic map(2, 5, 1)
    port map(
      index => fork5_outs_1,
      index_valid => fork5_outs_1_valid,
      index_ready => fork5_outs_1_ready,
      ins(0) => extsi52_outs,
      ins(1) => cond_br13_trueOut,
      ins_valid(0) => extsi52_outs_valid,
      ins_valid(1) => cond_br13_trueOut_valid,
      ins_ready(0) => extsi52_outs_ready,
      ins_ready(1) => cond_br13_trueOut_ready,
      clk => clk,
      rst => rst,
      outs => mux1_outs,
      outs_valid => mux1_outs_valid,
      outs_ready => mux1_outs_ready
    );

  buffer11 : entity work.tehb(arch) generic map(5)
    port map(
      ins => mux1_outs,
      ins_valid => mux1_outs_valid,
      ins_ready => mux1_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer11_outs,
      outs_valid => buffer11_outs_valid,
      outs_ready => buffer11_outs_ready
    );

  fork2 : entity work.handshake_fork(arch) generic map(2, 5)
    port map(
      ins => buffer11_outs,
      ins_valid => buffer11_outs_valid,
      ins_ready => buffer11_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork2_outs_0,
      outs(1) => fork2_outs_1,
      outs_valid(0) => fork2_outs_0_valid,
      outs_valid(1) => fork2_outs_1_valid,
      outs_ready(0) => fork2_outs_0_ready,
      outs_ready(1) => fork2_outs_1_ready
    );

  extsi54 : entity work.extsi(arch) generic map(5, 7)
    port map(
      ins => fork2_outs_0,
      ins_valid => fork2_outs_0_valid,
      ins_ready => fork2_outs_0_ready,
      clk => clk,
      rst => rst,
      outs => extsi54_outs,
      outs_valid => extsi54_outs_valid,
      outs_ready => extsi54_outs_ready
    );

  mux2 : entity work.mux(arch) generic map(2, 5, 1)
    port map(
      index => fork5_outs_0,
      index_valid => fork5_outs_0_valid,
      index_ready => fork5_outs_0_ready,
      ins(0) => buffer8_outs,
      ins(1) => cond_br14_trueOut,
      ins_valid(0) => buffer8_outs_valid,
      ins_valid(1) => cond_br14_trueOut_valid,
      ins_ready(0) => buffer8_outs_ready,
      ins_ready(1) => cond_br14_trueOut_ready,
      clk => clk,
      rst => rst,
      outs => mux2_outs,
      outs_valid => mux2_outs_valid,
      outs_ready => mux2_outs_ready
    );

  buffer12 : entity work.oehb(arch) generic map(5)
    port map(
      ins => mux2_outs,
      ins_valid => mux2_outs_valid,
      ins_ready => mux2_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer12_outs,
      outs_valid => buffer12_outs_valid,
      outs_ready => buffer12_outs_ready
    );

  buffer13 : entity work.tehb(arch) generic map(5)
    port map(
      ins => buffer12_outs,
      ins_valid => buffer12_outs_valid,
      ins_ready => buffer12_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer13_outs,
      outs_valid => buffer13_outs_valid,
      outs_ready => buffer13_outs_ready
    );

  fork3 : entity work.handshake_fork(arch) generic map(2, 5)
    port map(
      ins => buffer13_outs,
      ins_valid => buffer13_outs_valid,
      ins_ready => buffer13_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork3_outs_0,
      outs(1) => fork3_outs_1,
      outs_valid(0) => fork3_outs_0_valid,
      outs_valid(1) => fork3_outs_1_valid,
      outs_ready(0) => fork3_outs_0_ready,
      outs_ready(1) => fork3_outs_1_ready
    );

  extsi55 : entity work.extsi(arch) generic map(5, 32)
    port map(
      ins => fork3_outs_1,
      ins_valid => fork3_outs_1_valid,
      ins_ready => fork3_outs_1_ready,
      clk => clk,
      rst => rst,
      outs => extsi55_outs,
      outs_valid => extsi55_outs_valid,
      outs_ready => extsi55_outs_ready
    );

  fork4 : entity work.handshake_fork(arch) generic map(2, 32)
    port map(
      ins => extsi55_outs,
      ins_valid => extsi55_outs_valid,
      ins_ready => extsi55_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork4_outs_0,
      outs(1) => fork4_outs_1,
      outs_valid(0) => fork4_outs_0_valid,
      outs_valid(1) => fork4_outs_1_valid,
      outs_ready(0) => fork4_outs_0_ready,
      outs_ready(1) => fork4_outs_1_ready
    );

  control_merge1 : entity work.control_merge_dataless(arch) generic map(2, 1)
    port map(
      ins_valid(0) => fork1_outs_1_valid,
      ins_valid(1) => cond_br15_trueOut_valid,
      ins_ready(0) => fork1_outs_1_ready,
      ins_ready(1) => cond_br15_trueOut_ready,
      clk => clk,
      rst => rst,
      outs_valid => control_merge1_outs_valid,
      outs_ready => control_merge1_outs_ready,
      index => control_merge1_index,
      index_valid => control_merge1_index_valid,
      index_ready => control_merge1_index_ready
    );

  fork5 : entity work.handshake_fork(arch) generic map(2, 1)
    port map(
      ins => control_merge1_index,
      ins_valid => control_merge1_index_valid,
      ins_ready => control_merge1_index_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork5_outs_0,
      outs(1) => fork5_outs_1,
      outs_valid(0) => fork5_outs_0_valid,
      outs_valid(1) => fork5_outs_1_valid,
      outs_ready(0) => fork5_outs_0_ready,
      outs_ready(1) => fork5_outs_1_ready
    );

  fork6 : entity work.fork_dataless(arch) generic map(3)
    port map(
      ins_valid => control_merge1_outs_valid,
      ins_ready => control_merge1_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid(0) => fork6_outs_0_valid,
      outs_valid(1) => fork6_outs_1_valid,
      outs_valid(2) => fork6_outs_2_valid,
      outs_ready(0) => fork6_outs_0_ready,
      outs_ready(1) => fork6_outs_1_ready,
      outs_ready(2) => fork6_outs_2_ready
    );

  constant47 : entity work.handshake_constant_1(arch) generic map(2)
    port map(
      ctrl_valid => fork6_outs_1_valid,
      ctrl_ready => fork6_outs_1_ready,
      clk => clk,
      rst => rst,
      outs => constant47_outs,
      outs_valid => constant47_outs_valid,
      outs_ready => constant47_outs_ready
    );

  extsi2 : entity work.extsi(arch) generic map(2, 32)
    port map(
      ins => constant47_outs,
      ins_valid => constant47_outs_valid,
      ins_ready => constant47_outs_ready,
      clk => clk,
      rst => rst,
      outs => extsi2_outs,
      outs_valid => extsi2_outs_valid,
      outs_ready => extsi2_outs_ready
    );

  constant48 : entity work.handshake_constant_0(arch) generic map(1)
    port map(
      ctrl_valid => fork6_outs_0_valid,
      ctrl_ready => fork6_outs_0_ready,
      clk => clk,
      rst => rst,
      outs => constant48_outs,
      outs_valid => constant48_outs_valid,
      outs_ready => constant48_outs_ready
    );

  fork7 : entity work.handshake_fork(arch) generic map(2, 1)
    port map(
      ins => constant48_outs,
      ins_valid => constant48_outs_valid,
      ins_ready => constant48_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork7_outs_0,
      outs(1) => fork7_outs_1,
      outs_valid(0) => fork7_outs_0_valid,
      outs_valid(1) => fork7_outs_1_valid,
      outs_ready(0) => fork7_outs_0_ready,
      outs_ready(1) => fork7_outs_1_ready
    );

  extsi4 : entity work.extsi(arch) generic map(1, 32)
    port map(
      ins => fork7_outs_1,
      ins_valid => fork7_outs_1_valid,
      ins_ready => fork7_outs_1_ready,
      clk => clk,
      rst => rst,
      outs => extsi4_outs,
      outs_valid => extsi4_outs_valid,
      outs_ready => extsi4_outs_ready
    );

  source0 : entity work.source(arch)
    port map(
      clk => clk,
      rst => rst,
      outs_valid => source0_outs_valid,
      outs_ready => source0_outs_ready
    );

  constant49 : entity work.handshake_constant_1(arch) generic map(2)
    port map(
      ctrl_valid => source0_outs_valid,
      ctrl_ready => source0_outs_ready,
      clk => clk,
      rst => rst,
      outs => constant49_outs,
      outs_valid => constant49_outs_valid,
      outs_ready => constant49_outs_ready
    );

  extsi5 : entity work.extsi(arch) generic map(2, 32)
    port map(
      ins => constant49_outs,
      ins_valid => constant49_outs_valid,
      ins_ready => constant49_outs_ready,
      clk => clk,
      rst => rst,
      outs => extsi5_outs,
      outs_valid => extsi5_outs_valid,
      outs_ready => extsi5_outs_ready
    );

  source1 : entity work.source(arch)
    port map(
      clk => clk,
      rst => rst,
      outs_valid => source1_outs_valid,
      outs_ready => source1_outs_ready
    );

  constant50 : entity work.handshake_constant_2(arch) generic map(3)
    port map(
      ctrl_valid => source1_outs_valid,
      ctrl_ready => source1_outs_ready,
      clk => clk,
      rst => rst,
      outs => constant50_outs,
      outs_valid => constant50_outs_valid,
      outs_ready => constant50_outs_ready
    );

  extsi6 : entity work.extsi(arch) generic map(3, 32)
    port map(
      ins => constant50_outs,
      ins_valid => constant50_outs_valid,
      ins_ready => constant50_outs_ready,
      clk => clk,
      rst => rst,
      outs => extsi6_outs,
      outs_valid => extsi6_outs_valid,
      outs_ready => extsi6_outs_ready
    );

  shli0 : entity work.shli(arch) generic map(32)
    port map(
      lhs => fork4_outs_0,
      lhs_valid => fork4_outs_0_valid,
      lhs_ready => fork4_outs_0_ready,
      rhs => extsi5_outs,
      rhs_valid => extsi5_outs_valid,
      rhs_ready => extsi5_outs_ready,
      clk => clk,
      rst => rst,
      result => shli0_result,
      result_valid => shli0_result_valid,
      result_ready => shli0_result_ready
    );

  buffer14 : entity work.oehb(arch) generic map(32)
    port map(
      ins => shli0_result,
      ins_valid => shli0_result_valid,
      ins_ready => shli0_result_ready,
      clk => clk,
      rst => rst,
      outs => buffer14_outs,
      outs_valid => buffer14_outs_valid,
      outs_ready => buffer14_outs_ready
    );

  trunci0 : entity work.trunci(arch) generic map(32, 7)
    port map(
      ins => buffer14_outs,
      ins_valid => buffer14_outs_valid,
      ins_ready => buffer14_outs_ready,
      clk => clk,
      rst => rst,
      outs => trunci0_outs,
      outs_valid => trunci0_outs_valid,
      outs_ready => trunci0_outs_ready
    );

  shli1 : entity work.shli(arch) generic map(32)
    port map(
      lhs => fork4_outs_1,
      lhs_valid => fork4_outs_1_valid,
      lhs_ready => fork4_outs_1_ready,
      rhs => extsi6_outs,
      rhs_valid => extsi6_outs_valid,
      rhs_ready => extsi6_outs_ready,
      clk => clk,
      rst => rst,
      result => shli1_result,
      result_valid => shli1_result_valid,
      result_ready => shli1_result_ready
    );

  buffer15 : entity work.oehb(arch) generic map(32)
    port map(
      ins => shli1_result,
      ins_valid => shli1_result_valid,
      ins_ready => shli1_result_ready,
      clk => clk,
      rst => rst,
      outs => buffer15_outs,
      outs_valid => buffer15_outs_valid,
      outs_ready => buffer15_outs_ready
    );

  trunci1 : entity work.trunci(arch) generic map(32, 7)
    port map(
      ins => buffer15_outs,
      ins_valid => buffer15_outs_valid,
      ins_ready => buffer15_outs_ready,
      clk => clk,
      rst => rst,
      outs => trunci1_outs,
      outs_valid => trunci1_outs_valid,
      outs_ready => trunci1_outs_ready
    );

  addi27 : entity work.addi(arch) generic map(7)
    port map(
      lhs => trunci0_outs,
      lhs_valid => trunci0_outs_valid,
      lhs_ready => trunci0_outs_ready,
      rhs => trunci1_outs,
      rhs_valid => trunci1_outs_valid,
      rhs_ready => trunci1_outs_ready,
      clk => clk,
      rst => rst,
      result => addi27_result,
      result_valid => addi27_result_valid,
      result_ready => addi27_result_ready
    );

  buffer16 : entity work.oehb(arch) generic map(7)
    port map(
      ins => addi27_result,
      ins_valid => addi27_result_valid,
      ins_ready => addi27_result_ready,
      clk => clk,
      rst => rst,
      outs => buffer16_outs,
      outs_valid => buffer16_outs_valid,
      outs_ready => buffer16_outs_ready
    );

  addi3 : entity work.addi(arch) generic map(7)
    port map(
      lhs => extsi54_outs,
      lhs_valid => extsi54_outs_valid,
      lhs_ready => extsi54_outs_ready,
      rhs => buffer16_outs,
      rhs_valid => buffer16_outs_valid,
      rhs_ready => buffer16_outs_ready,
      clk => clk,
      rst => rst,
      result => addi3_result,
      result_valid => addi3_result_valid,
      result_ready => addi3_result_ready
    );

  buffer0 : entity work.tfifo_dataless(arch) generic map(1)
    port map(
      ins_valid => store0_doneOut_valid,
      ins_ready => store0_doneOut_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer0_outs_valid,
      outs_ready => buffer0_outs_ready
    );

  fork8 : entity work.fork_dataless(arch) generic map(2)
    port map(
      ins_valid => buffer0_outs_valid,
      ins_ready => buffer0_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid(0) => fork8_outs_0_valid,
      outs_valid(1) => fork8_outs_1_valid,
      outs_ready(0) => fork8_outs_0_ready,
      outs_ready(1) => fork8_outs_1_ready
    );

  buffer17 : entity work.oehb(arch) generic map(7)
    port map(
      ins => addi3_result,
      ins_valid => addi3_result_valid,
      ins_ready => addi3_result_ready,
      clk => clk,
      rst => rst,
      outs => buffer17_outs,
      outs_valid => buffer17_outs_valid,
      outs_ready => buffer17_outs_ready
    );

  store0 : entity work.store(arch) generic map(32, 7)
    port map(
      addrIn => buffer17_outs,
      addrIn_valid => buffer17_outs_valid,
      addrIn_ready => buffer17_outs_ready,
      dataIn => extsi4_outs,
      dataIn_valid => extsi4_outs_valid,
      dataIn_ready => extsi4_outs_ready,
      doneFromMem_valid => mem_controller6_stDone_0_valid,
      doneFromMem_ready => mem_controller6_stDone_0_ready,
      clk => clk,
      rst => rst,
      addrOut => store0_addrOut,
      addrOut_valid => store0_addrOut_valid,
      addrOut_ready => store0_addrOut_ready,
      dataToMem => store0_dataToMem,
      dataToMem_valid => store0_dataToMem_valid,
      dataToMem_ready => store0_dataToMem_ready,
      doneOut_valid => store0_doneOut_valid,
      doneOut_ready => store0_doneOut_ready
    );

  extsi51 : entity work.extsi(arch) generic map(1, 5)
    port map(
      ins => fork7_outs_0,
      ins_valid => fork7_outs_0_valid,
      ins_ready => fork7_outs_0_ready,
      clk => clk,
      rst => rst,
      outs => extsi51_outs,
      outs_valid => extsi51_outs_valid,
      outs_ready => extsi51_outs_ready
    );

  buffer65 : entity work.oehb_dataless(arch)
    port map(
      ins_valid => buffer1_outs_valid,
      ins_ready => buffer1_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer65_outs_valid,
      outs_ready => buffer65_outs_ready
    );

  cond_br116 : entity work.cond_br_dataless(arch)
    port map(
      condition => buffer18_outs,
      condition_valid => buffer18_outs_valid,
      condition_ready => buffer18_outs_ready,
      data_valid => buffer65_outs_valid,
      data_ready => buffer65_outs_ready,
      clk => clk,
      rst => rst,
      trueOut_valid => cond_br116_trueOut_valid,
      trueOut_ready => cond_br116_trueOut_ready,
      falseOut_valid => cond_br116_falseOut_valid,
      falseOut_ready => cond_br116_falseOut_ready
    );

  buffer18 : entity work.tfifo(arch) generic map(4, 1)
    port map(
      ins => fork23_outs_5,
      ins_valid => fork23_outs_5_valid,
      ins_ready => fork23_outs_5_ready,
      clk => clk,
      rst => rst,
      outs => buffer18_outs,
      outs_valid => buffer18_outs_valid,
      outs_ready => buffer18_outs_ready
    );

  cond_br117 : entity work.cond_br_dataless(arch)
    port map(
      condition => buffer19_outs,
      condition_valid => buffer19_outs_valid,
      condition_ready => buffer19_outs_ready,
      data_valid => fork10_outs_2_valid,
      data_ready => fork10_outs_2_ready,
      clk => clk,
      rst => rst,
      trueOut_valid => cond_br117_trueOut_valid,
      trueOut_ready => cond_br117_trueOut_ready,
      falseOut_valid => cond_br117_falseOut_valid,
      falseOut_ready => cond_br117_falseOut_ready
    );

  buffer19 : entity work.tfifo(arch) generic map(3, 1)
    port map(
      ins => fork23_outs_4,
      ins_valid => fork23_outs_4_valid,
      ins_ready => fork23_outs_4_ready,
      clk => clk,
      rst => rst,
      outs => buffer19_outs,
      outs_valid => buffer19_outs_valid,
      outs_ready => buffer19_outs_ready
    );

  sink0 : entity work.sink_dataless(arch)
    port map(
      ins_valid => cond_br117_falseOut_valid,
      ins_ready => cond_br117_falseOut_ready,
      clk => clk,
      rst => rst
    );

  init10 : entity work.tehb_init(arch) generic map(1, 0)
    port map(
      ins => fork23_outs_3,
      ins_valid => fork23_outs_3_valid,
      ins_ready => fork23_outs_3_ready,
      clk => clk,
      rst => rst,
      outs => init10_outs,
      outs_valid => init10_outs_valid,
      outs_ready => init10_outs_ready
    );

  fork9 : entity work.handshake_fork(arch) generic map(2, 1)
    port map(
      ins => init10_outs,
      ins_valid => init10_outs_valid,
      ins_ready => init10_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork9_outs_0,
      outs(1) => fork9_outs_1,
      outs_valid(0) => fork9_outs_0_valid,
      outs_valid(1) => fork9_outs_1_valid,
      outs_ready(0) => fork9_outs_0_ready,
      outs_ready(1) => fork9_outs_1_ready
    );

  mux28 : entity work.mux_dataless(arch) generic map(2, 1)
    port map(
      index => buffer21_outs,
      index_valid => buffer21_outs_valid,
      index_ready => buffer21_outs_ready,
      ins_valid(0) => fork8_outs_1_valid,
      ins_valid(1) => cond_br117_trueOut_valid,
      ins_ready(0) => fork8_outs_1_ready,
      ins_ready(1) => cond_br117_trueOut_ready,
      clk => clk,
      rst => rst,
      outs_valid => mux28_outs_valid,
      outs_ready => mux28_outs_ready
    );

  buffer21 : entity work.tfifo(arch) generic map(3, 1)
    port map(
      ins => fork9_outs_1,
      ins_valid => fork9_outs_1_valid,
      ins_ready => fork9_outs_1_ready,
      clk => clk,
      rst => rst,
      outs => buffer21_outs,
      outs_valid => buffer21_outs_valid,
      outs_ready => buffer21_outs_ready
    );

  buffer20 : entity work.oehb_dataless(arch)
    port map(
      ins_valid => mux28_outs_valid,
      ins_ready => mux28_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer20_outs_valid,
      outs_ready => buffer20_outs_ready
    );

  buffer23 : entity work.tehb_dataless(arch)
    port map(
      ins_valid => buffer20_outs_valid,
      ins_ready => buffer20_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer23_outs_valid,
      outs_ready => buffer23_outs_ready
    );

  fork10 : entity work.fork_dataless(arch) generic map(3)
    port map(
      ins_valid => buffer23_outs_valid,
      ins_ready => buffer23_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid(0) => fork10_outs_0_valid,
      outs_valid(1) => fork10_outs_1_valid,
      outs_valid(2) => fork10_outs_2_valid,
      outs_ready(0) => fork10_outs_0_ready,
      outs_ready(1) => fork10_outs_1_ready,
      outs_ready(2) => fork10_outs_2_ready
    );

  buffer9 : entity work.oehb_dataless(arch)
    port map(
      ins_valid => mux27_outs_valid,
      ins_ready => mux27_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer9_outs_valid,
      outs_ready => buffer9_outs_ready
    );

  buffer10 : entity work.tehb_dataless(arch)
    port map(
      ins_valid => buffer9_outs_valid,
      ins_ready => buffer9_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer10_outs_valid,
      outs_ready => buffer10_outs_ready
    );

  mux31 : entity work.mux_dataless(arch) generic map(2, 1)
    port map(
      index => buffer22_outs,
      index_valid => buffer22_outs_valid,
      index_ready => buffer22_outs_ready,
      ins_valid(0) => buffer10_outs_valid,
      ins_valid(1) => cond_br116_trueOut_valid,
      ins_ready(0) => buffer10_outs_ready,
      ins_ready(1) => cond_br116_trueOut_ready,
      clk => clk,
      rst => rst,
      outs_valid => mux31_outs_valid,
      outs_ready => mux31_outs_ready
    );

  buffer22 : entity work.tfifo(arch) generic map(4, 1)
    port map(
      ins => fork9_outs_0,
      ins_valid => fork9_outs_0_valid,
      ins_ready => fork9_outs_0_ready,
      clk => clk,
      rst => rst,
      outs => buffer22_outs,
      outs_valid => buffer22_outs_valid,
      outs_ready => buffer22_outs_ready
    );

  mux3 : entity work.mux(arch) generic map(2, 5, 1)
    port map(
      index => fork17_outs_2,
      index_valid => fork17_outs_2_valid,
      index_ready => fork17_outs_2_ready,
      ins(0) => extsi51_outs,
      ins(1) => cond_br9_trueOut,
      ins_valid(0) => extsi51_outs_valid,
      ins_valid(1) => cond_br9_trueOut_valid,
      ins_ready(0) => extsi51_outs_ready,
      ins_ready(1) => cond_br9_trueOut_ready,
      clk => clk,
      rst => rst,
      outs => mux3_outs,
      outs_valid => mux3_outs_valid,
      outs_ready => mux3_outs_ready
    );

  buffer26 : entity work.oehb(arch) generic map(5)
    port map(
      ins => mux3_outs,
      ins_valid => mux3_outs_valid,
      ins_ready => mux3_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer26_outs,
      outs_valid => buffer26_outs_valid,
      outs_ready => buffer26_outs_ready
    );

  buffer27 : entity work.tehb(arch) generic map(5)
    port map(
      ins => buffer26_outs,
      ins_valid => buffer26_outs_valid,
      ins_ready => buffer26_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer27_outs,
      outs_valid => buffer27_outs_valid,
      outs_ready => buffer27_outs_ready
    );

  fork11 : entity work.handshake_fork(arch) generic map(3, 5)
    port map(
      ins => buffer27_outs,
      ins_valid => buffer27_outs_valid,
      ins_ready => buffer27_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork11_outs_0,
      outs(1) => fork11_outs_1,
      outs(2) => fork11_outs_2,
      outs_valid(0) => fork11_outs_0_valid,
      outs_valid(1) => fork11_outs_1_valid,
      outs_valid(2) => fork11_outs_2_valid,
      outs_ready(0) => fork11_outs_0_ready,
      outs_ready(1) => fork11_outs_1_ready,
      outs_ready(2) => fork11_outs_2_ready
    );

  extsi56 : entity work.extsi(arch) generic map(5, 7)
    port map(
      ins => buffer24_outs,
      ins_valid => buffer24_outs_valid,
      ins_ready => buffer24_outs_ready,
      clk => clk,
      rst => rst,
      outs => extsi56_outs,
      outs_valid => extsi56_outs_valid,
      outs_ready => extsi56_outs_ready
    );

  buffer24 : entity work.tfifo(arch) generic map(1, 5)
    port map(
      ins => fork11_outs_0,
      ins_valid => fork11_outs_0_valid,
      ins_ready => fork11_outs_0_ready,
      clk => clk,
      rst => rst,
      outs => buffer24_outs,
      outs_valid => buffer24_outs_valid,
      outs_ready => buffer24_outs_ready
    );

  extsi57 : entity work.extsi(arch) generic map(5, 6)
    port map(
      ins => fork11_outs_1,
      ins_valid => fork11_outs_1_valid,
      ins_ready => fork11_outs_1_ready,
      clk => clk,
      rst => rst,
      outs => extsi57_outs,
      outs_valid => extsi57_outs_valid,
      outs_ready => extsi57_outs_ready
    );

  extsi58 : entity work.extsi(arch) generic map(5, 32)
    port map(
      ins => fork11_outs_2,
      ins_valid => fork11_outs_2_valid,
      ins_ready => fork11_outs_2_ready,
      clk => clk,
      rst => rst,
      outs => extsi58_outs,
      outs_valid => extsi58_outs_valid,
      outs_ready => extsi58_outs_ready
    );

  fork12 : entity work.handshake_fork(arch) generic map(2, 32)
    port map(
      ins => extsi58_outs,
      ins_valid => extsi58_outs_valid,
      ins_ready => extsi58_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork12_outs_0,
      outs(1) => fork12_outs_1,
      outs_valid(0) => fork12_outs_0_valid,
      outs_valid(1) => fork12_outs_1_valid,
      outs_ready(0) => fork12_outs_0_ready,
      outs_ready(1) => fork12_outs_1_ready
    );

  mux4 : entity work.mux(arch) generic map(2, 5, 1)
    port map(
      index => fork17_outs_0,
      index_valid => fork17_outs_0_valid,
      index_ready => fork17_outs_0_ready,
      ins(0) => fork3_outs_0,
      ins(1) => cond_br10_trueOut,
      ins_valid(0) => fork3_outs_0_valid,
      ins_valid(1) => cond_br10_trueOut_valid,
      ins_ready(0) => fork3_outs_0_ready,
      ins_ready(1) => cond_br10_trueOut_ready,
      clk => clk,
      rst => rst,
      outs => mux4_outs,
      outs_valid => mux4_outs_valid,
      outs_ready => mux4_outs_ready
    );

  buffer28 : entity work.oehb(arch) generic map(5)
    port map(
      ins => mux4_outs,
      ins_valid => mux4_outs_valid,
      ins_ready => mux4_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer28_outs,
      outs_valid => buffer28_outs_valid,
      outs_ready => buffer28_outs_ready
    );

  buffer29 : entity work.tehb(arch) generic map(5)
    port map(
      ins => buffer28_outs,
      ins_valid => buffer28_outs_valid,
      ins_ready => buffer28_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer29_outs,
      outs_valid => buffer29_outs_valid,
      outs_ready => buffer29_outs_ready
    );

  fork13 : entity work.handshake_fork(arch) generic map(2, 5)
    port map(
      ins => buffer29_outs,
      ins_valid => buffer29_outs_valid,
      ins_ready => buffer29_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork13_outs_0,
      outs(1) => fork13_outs_1,
      outs_valid(0) => fork13_outs_0_valid,
      outs_valid(1) => fork13_outs_1_valid,
      outs_ready(0) => fork13_outs_0_ready,
      outs_ready(1) => fork13_outs_1_ready
    );

  extsi59 : entity work.extsi(arch) generic map(5, 32)
    port map(
      ins => fork13_outs_1,
      ins_valid => fork13_outs_1_valid,
      ins_ready => fork13_outs_1_ready,
      clk => clk,
      rst => rst,
      outs => extsi59_outs,
      outs_valid => extsi59_outs_valid,
      outs_ready => extsi59_outs_ready
    );

  fork14 : entity work.handshake_fork(arch) generic map(6, 32)
    port map(
      ins => extsi59_outs,
      ins_valid => extsi59_outs_valid,
      ins_ready => extsi59_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork14_outs_0,
      outs(1) => fork14_outs_1,
      outs(2) => fork14_outs_2,
      outs(3) => fork14_outs_3,
      outs(4) => fork14_outs_4,
      outs(5) => fork14_outs_5,
      outs_valid(0) => fork14_outs_0_valid,
      outs_valid(1) => fork14_outs_1_valid,
      outs_valid(2) => fork14_outs_2_valid,
      outs_valid(3) => fork14_outs_3_valid,
      outs_valid(4) => fork14_outs_4_valid,
      outs_valid(5) => fork14_outs_5_valid,
      outs_ready(0) => fork14_outs_0_ready,
      outs_ready(1) => fork14_outs_1_ready,
      outs_ready(2) => fork14_outs_2_ready,
      outs_ready(3) => fork14_outs_3_ready,
      outs_ready(4) => fork14_outs_4_ready,
      outs_ready(5) => fork14_outs_5_ready
    );

  mux5 : entity work.mux(arch) generic map(2, 5, 1)
    port map(
      index => fork17_outs_1,
      index_valid => fork17_outs_1_valid,
      index_ready => fork17_outs_1_ready,
      ins(0) => fork2_outs_1,
      ins(1) => cond_br11_trueOut,
      ins_valid(0) => fork2_outs_1_valid,
      ins_valid(1) => cond_br11_trueOut_valid,
      ins_ready(0) => fork2_outs_1_ready,
      ins_ready(1) => cond_br11_trueOut_ready,
      clk => clk,
      rst => rst,
      outs => mux5_outs,
      outs_valid => mux5_outs_valid,
      outs_ready => mux5_outs_ready
    );

  buffer31 : entity work.oehb(arch) generic map(5)
    port map(
      ins => mux5_outs,
      ins_valid => mux5_outs_valid,
      ins_ready => mux5_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer31_outs,
      outs_valid => buffer31_outs_valid,
      outs_ready => buffer31_outs_ready
    );

  buffer34 : entity work.tehb(arch) generic map(5)
    port map(
      ins => buffer31_outs,
      ins_valid => buffer31_outs_valid,
      ins_ready => buffer31_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer34_outs,
      outs_valid => buffer34_outs_valid,
      outs_ready => buffer34_outs_ready
    );

  fork15 : entity work.handshake_fork(arch) generic map(3, 5)
    port map(
      ins => buffer34_outs,
      ins_valid => buffer34_outs_valid,
      ins_ready => buffer34_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork15_outs_0,
      outs(1) => fork15_outs_1,
      outs(2) => fork15_outs_2,
      outs_valid(0) => fork15_outs_0_valid,
      outs_valid(1) => fork15_outs_1_valid,
      outs_valid(2) => fork15_outs_2_valid,
      outs_ready(0) => fork15_outs_0_ready,
      outs_ready(1) => fork15_outs_1_ready,
      outs_ready(2) => fork15_outs_2_ready
    );

  extsi60 : entity work.extsi(arch) generic map(5, 7)
    port map(
      ins => buffer30_outs,
      ins_valid => buffer30_outs_valid,
      ins_ready => buffer30_outs_ready,
      clk => clk,
      rst => rst,
      outs => extsi60_outs,
      outs_valid => extsi60_outs_valid,
      outs_ready => extsi60_outs_ready
    );

  buffer30 : entity work.tfifo(arch) generic map(1, 5)
    port map(
      ins => fork15_outs_0,
      ins_valid => fork15_outs_0_valid,
      ins_ready => fork15_outs_0_ready,
      clk => clk,
      rst => rst,
      outs => buffer30_outs,
      outs_valid => buffer30_outs_valid,
      outs_ready => buffer30_outs_ready
    );

  extsi61 : entity work.extsi(arch) generic map(5, 32)
    port map(
      ins => fork15_outs_2,
      ins_valid => fork15_outs_2_valid,
      ins_ready => fork15_outs_2_ready,
      clk => clk,
      rst => rst,
      outs => extsi61_outs,
      outs_valid => extsi61_outs_valid,
      outs_ready => extsi61_outs_ready
    );

  fork16 : entity work.handshake_fork(arch) generic map(2, 32)
    port map(
      ins => extsi61_outs,
      ins_valid => extsi61_outs_valid,
      ins_ready => extsi61_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork16_outs_0,
      outs(1) => fork16_outs_1,
      outs_valid(0) => fork16_outs_0_valid,
      outs_valid(1) => fork16_outs_1_valid,
      outs_ready(0) => fork16_outs_0_ready,
      outs_ready(1) => fork16_outs_1_ready
    );

  control_merge2 : entity work.control_merge_dataless(arch) generic map(2, 1)
    port map(
      ins_valid(0) => fork6_outs_2_valid,
      ins_valid(1) => cond_br12_trueOut_valid,
      ins_ready(0) => fork6_outs_2_ready,
      ins_ready(1) => cond_br12_trueOut_ready,
      clk => clk,
      rst => rst,
      outs_valid => control_merge2_outs_valid,
      outs_ready => control_merge2_outs_ready,
      index => control_merge2_index,
      index_valid => control_merge2_index_valid,
      index_ready => control_merge2_index_ready
    );

  fork17 : entity work.handshake_fork(arch) generic map(3, 1)
    port map(
      ins => control_merge2_index,
      ins_valid => control_merge2_index_valid,
      ins_ready => control_merge2_index_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork17_outs_0,
      outs(1) => fork17_outs_1,
      outs(2) => fork17_outs_2,
      outs_valid(0) => fork17_outs_0_valid,
      outs_valid(1) => fork17_outs_1_valid,
      outs_valid(2) => fork17_outs_2_valid,
      outs_ready(0) => fork17_outs_0_ready,
      outs_ready(1) => fork17_outs_1_ready,
      outs_ready(2) => fork17_outs_2_ready
    );

  fork18 : entity work.fork_dataless(arch) generic map(2)
    port map(
      ins_valid => control_merge2_outs_valid,
      ins_ready => control_merge2_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid(0) => fork18_outs_0_valid,
      outs_valid(1) => fork18_outs_1_valid,
      outs_ready(0) => fork18_outs_0_ready,
      outs_ready(1) => fork18_outs_1_ready
    );

  constant51 : entity work.handshake_constant_1(arch) generic map(2)
    port map(
      ctrl_valid => fork18_outs_0_valid,
      ctrl_ready => fork18_outs_0_ready,
      clk => clk,
      rst => rst,
      outs => constant51_outs,
      outs_valid => constant51_outs_valid,
      outs_ready => constant51_outs_ready
    );

  extsi7 : entity work.extsi(arch) generic map(2, 32)
    port map(
      ins => constant51_outs,
      ins_valid => constant51_outs_valid,
      ins_ready => constant51_outs_ready,
      clk => clk,
      rst => rst,
      outs => extsi7_outs,
      outs_valid => extsi7_outs_valid,
      outs_ready => extsi7_outs_ready
    );

  source2 : entity work.source(arch)
    port map(
      clk => clk,
      rst => rst,
      outs_valid => source2_outs_valid,
      outs_ready => source2_outs_ready
    );

  constant52 : entity work.handshake_constant_3(arch) generic map(5)
    port map(
      ctrl_valid => source2_outs_valid,
      ctrl_ready => source2_outs_ready,
      clk => clk,
      rst => rst,
      outs => constant52_outs,
      outs_valid => constant52_outs_valid,
      outs_ready => constant52_outs_ready
    );

  extsi62 : entity work.extsi(arch) generic map(5, 6)
    port map(
      ins => constant52_outs,
      ins_valid => constant52_outs_valid,
      ins_ready => constant52_outs_ready,
      clk => clk,
      rst => rst,
      outs => extsi62_outs,
      outs_valid => extsi62_outs_valid,
      outs_ready => extsi62_outs_ready
    );

  source3 : entity work.source(arch)
    port map(
      clk => clk,
      rst => rst,
      outs_valid => source3_outs_valid,
      outs_ready => source3_outs_ready
    );

  constant53 : entity work.handshake_constant_1(arch) generic map(2)
    port map(
      ctrl_valid => source3_outs_valid,
      ctrl_ready => source3_outs_ready,
      clk => clk,
      rst => rst,
      outs => constant53_outs,
      outs_valid => constant53_outs_valid,
      outs_ready => constant53_outs_ready
    );

  fork19 : entity work.handshake_fork(arch) generic map(2, 2)
    port map(
      ins => constant53_outs,
      ins_valid => constant53_outs_valid,
      ins_ready => constant53_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork19_outs_0,
      outs(1) => fork19_outs_1,
      outs_valid(0) => fork19_outs_0_valid,
      outs_valid(1) => fork19_outs_1_valid,
      outs_ready(0) => fork19_outs_0_ready,
      outs_ready(1) => fork19_outs_1_ready
    );

  extsi63 : entity work.extsi(arch) generic map(2, 6)
    port map(
      ins => buffer32_outs,
      ins_valid => buffer32_outs_valid,
      ins_ready => buffer32_outs_ready,
      clk => clk,
      rst => rst,
      outs => extsi63_outs,
      outs_valid => extsi63_outs_valid,
      outs_ready => extsi63_outs_ready
    );

  buffer32 : entity work.tfifo(arch) generic map(1, 2)
    port map(
      ins => fork19_outs_0,
      ins_valid => fork19_outs_0_valid,
      ins_ready => fork19_outs_0_ready,
      clk => clk,
      rst => rst,
      outs => buffer32_outs,
      outs_valid => buffer32_outs_valid,
      outs_ready => buffer32_outs_ready
    );

  extsi9 : entity work.extsi(arch) generic map(2, 32)
    port map(
      ins => buffer33_outs,
      ins_valid => buffer33_outs_valid,
      ins_ready => buffer33_outs_ready,
      clk => clk,
      rst => rst,
      outs => extsi9_outs,
      outs_valid => extsi9_outs_valid,
      outs_ready => extsi9_outs_ready
    );

  buffer33 : entity work.tfifo(arch) generic map(1, 2)
    port map(
      ins => fork19_outs_1,
      ins_valid => fork19_outs_1_valid,
      ins_ready => fork19_outs_1_ready,
      clk => clk,
      rst => rst,
      outs => buffer33_outs,
      outs_valid => buffer33_outs_valid,
      outs_ready => buffer33_outs_ready
    );

  fork20 : entity work.handshake_fork(arch) generic map(4, 32)
    port map(
      ins => extsi9_outs,
      ins_valid => extsi9_outs_valid,
      ins_ready => extsi9_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork20_outs_0,
      outs(1) => fork20_outs_1,
      outs(2) => fork20_outs_2,
      outs(3) => fork20_outs_3,
      outs_valid(0) => fork20_outs_0_valid,
      outs_valid(1) => fork20_outs_1_valid,
      outs_valid(2) => fork20_outs_2_valid,
      outs_valid(3) => fork20_outs_3_valid,
      outs_ready(0) => fork20_outs_0_ready,
      outs_ready(1) => fork20_outs_1_ready,
      outs_ready(2) => fork20_outs_2_ready,
      outs_ready(3) => fork20_outs_3_ready
    );

  source4 : entity work.source(arch)
    port map(
      clk => clk,
      rst => rst,
      outs_valid => source4_outs_valid,
      outs_ready => source4_outs_ready
    );

  constant54 : entity work.handshake_constant_2(arch) generic map(3)
    port map(
      ctrl_valid => source4_outs_valid,
      ctrl_ready => source4_outs_ready,
      clk => clk,
      rst => rst,
      outs => constant54_outs,
      outs_valid => constant54_outs_valid,
      outs_ready => constant54_outs_ready
    );

  extsi10 : entity work.extsi(arch) generic map(3, 32)
    port map(
      ins => constant54_outs,
      ins_valid => constant54_outs_valid,
      ins_ready => constant54_outs_ready,
      clk => clk,
      rst => rst,
      outs => extsi10_outs,
      outs_valid => extsi10_outs_valid,
      outs_ready => extsi10_outs_ready
    );

  fork21 : entity work.handshake_fork(arch) generic map(4, 32)
    port map(
      ins => extsi10_outs,
      ins_valid => extsi10_outs_valid,
      ins_ready => extsi10_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork21_outs_0,
      outs(1) => fork21_outs_1,
      outs(2) => fork21_outs_2,
      outs(3) => fork21_outs_3,
      outs_valid(0) => fork21_outs_0_valid,
      outs_valid(1) => fork21_outs_1_valid,
      outs_valid(2) => fork21_outs_2_valid,
      outs_valid(3) => fork21_outs_3_valid,
      outs_ready(0) => fork21_outs_0_ready,
      outs_ready(1) => fork21_outs_1_ready,
      outs_ready(2) => fork21_outs_2_ready,
      outs_ready(3) => fork21_outs_3_ready
    );

  shli2 : entity work.shli(arch) generic map(32)
    port map(
      lhs => buffer35_outs,
      lhs_valid => buffer35_outs_valid,
      lhs_ready => buffer35_outs_ready,
      rhs => fork20_outs_0,
      rhs_valid => fork20_outs_0_valid,
      rhs_ready => fork20_outs_0_ready,
      clk => clk,
      rst => rst,
      result => shli2_result,
      result_valid => shli2_result_valid,
      result_ready => shli2_result_ready
    );

  buffer35 : entity work.tfifo(arch) generic map(1, 32)
    port map(
      ins => fork14_outs_0,
      ins_valid => fork14_outs_0_valid,
      ins_ready => fork14_outs_0_ready,
      clk => clk,
      rst => rst,
      outs => buffer35_outs,
      outs_valid => buffer35_outs_valid,
      outs_ready => buffer35_outs_ready
    );

  buffer38 : entity work.oehb(arch) generic map(32)
    port map(
      ins => shli2_result,
      ins_valid => shli2_result_valid,
      ins_ready => shli2_result_ready,
      clk => clk,
      rst => rst,
      outs => buffer38_outs,
      outs_valid => buffer38_outs_valid,
      outs_ready => buffer38_outs_ready
    );

  trunci2 : entity work.trunci(arch) generic map(32, 7)
    port map(
      ins => buffer38_outs,
      ins_valid => buffer38_outs_valid,
      ins_ready => buffer38_outs_ready,
      clk => clk,
      rst => rst,
      outs => trunci2_outs,
      outs_valid => trunci2_outs_valid,
      outs_ready => trunci2_outs_ready
    );

  shli3 : entity work.shli(arch) generic map(32)
    port map(
      lhs => buffer37_outs,
      lhs_valid => buffer37_outs_valid,
      lhs_ready => buffer37_outs_ready,
      rhs => fork21_outs_0,
      rhs_valid => fork21_outs_0_valid,
      rhs_ready => fork21_outs_0_ready,
      clk => clk,
      rst => rst,
      result => shli3_result,
      result_valid => shli3_result_valid,
      result_ready => shli3_result_ready
    );

  buffer37 : entity work.tfifo(arch) generic map(1, 32)
    port map(
      ins => fork14_outs_1,
      ins_valid => fork14_outs_1_valid,
      ins_ready => fork14_outs_1_ready,
      clk => clk,
      rst => rst,
      outs => buffer37_outs,
      outs_valid => buffer37_outs_valid,
      outs_ready => buffer37_outs_ready
    );

  buffer40 : entity work.oehb(arch) generic map(32)
    port map(
      ins => shli3_result,
      ins_valid => shli3_result_valid,
      ins_ready => shli3_result_ready,
      clk => clk,
      rst => rst,
      outs => buffer40_outs,
      outs_valid => buffer40_outs_valid,
      outs_ready => buffer40_outs_ready
    );

  trunci3 : entity work.trunci(arch) generic map(32, 7)
    port map(
      ins => buffer40_outs,
      ins_valid => buffer40_outs_valid,
      ins_ready => buffer40_outs_ready,
      clk => clk,
      rst => rst,
      outs => trunci3_outs,
      outs_valid => trunci3_outs_valid,
      outs_ready => trunci3_outs_ready
    );

  addi28 : entity work.addi(arch) generic map(7)
    port map(
      lhs => trunci2_outs,
      lhs_valid => trunci2_outs_valid,
      lhs_ready => trunci2_outs_ready,
      rhs => trunci3_outs,
      rhs_valid => trunci3_outs_valid,
      rhs_ready => trunci3_outs_ready,
      clk => clk,
      rst => rst,
      result => addi28_result,
      result_valid => addi28_result_valid,
      result_ready => addi28_result_ready
    );

  buffer52 : entity work.oehb(arch) generic map(7)
    port map(
      ins => addi28_result,
      ins_valid => addi28_result_valid,
      ins_ready => addi28_result_ready,
      clk => clk,
      rst => rst,
      outs => buffer52_outs,
      outs_valid => buffer52_outs_valid,
      outs_ready => buffer52_outs_ready
    );

  addi4 : entity work.addi(arch) generic map(7)
    port map(
      lhs => extsi56_outs,
      lhs_valid => extsi56_outs_valid,
      lhs_ready => extsi56_outs_ready,
      rhs => buffer52_outs,
      rhs_valid => buffer52_outs_valid,
      rhs_ready => buffer52_outs_ready,
      clk => clk,
      rst => rst,
      result => addi4_result,
      result_valid => addi4_result_valid,
      result_ready => addi4_result_ready
    );

  load0 : entity work.load(arch) generic map(32, 7)
    port map(
      addrIn => addi4_result,
      addrIn_valid => addi4_result_valid,
      addrIn_ready => addi4_result_ready,
      dataFromMem => mem_controller10_ldData_0,
      dataFromMem_valid => mem_controller10_ldData_0_valid,
      dataFromMem_ready => mem_controller10_ldData_0_ready,
      clk => clk,
      rst => rst,
      addrOut => load0_addrOut,
      addrOut_valid => load0_addrOut_valid,
      addrOut_ready => load0_addrOut_ready,
      dataOut => load0_dataOut,
      dataOut_valid => load0_dataOut_valid,
      dataOut_ready => load0_dataOut_ready
    );

  shli4 : entity work.shli(arch) generic map(32)
    port map(
      lhs => buffer39_outs,
      lhs_valid => buffer39_outs_valid,
      lhs_ready => buffer39_outs_ready,
      rhs => fork20_outs_1,
      rhs_valid => fork20_outs_1_valid,
      rhs_ready => fork20_outs_1_ready,
      clk => clk,
      rst => rst,
      result => shli4_result,
      result_valid => shli4_result_valid,
      result_ready => shli4_result_ready
    );

  buffer39 : entity work.tfifo(arch) generic map(1, 32)
    port map(
      ins => fork12_outs_0,
      ins_valid => fork12_outs_0_valid,
      ins_ready => fork12_outs_0_ready,
      clk => clk,
      rst => rst,
      outs => buffer39_outs,
      outs_valid => buffer39_outs_valid,
      outs_ready => buffer39_outs_ready
    );

  buffer53 : entity work.oehb(arch) generic map(32)
    port map(
      ins => shli4_result,
      ins_valid => shli4_result_valid,
      ins_ready => shli4_result_ready,
      clk => clk,
      rst => rst,
      outs => buffer53_outs,
      outs_valid => buffer53_outs_valid,
      outs_ready => buffer53_outs_ready
    );

  trunci4 : entity work.trunci(arch) generic map(32, 7)
    port map(
      ins => buffer53_outs,
      ins_valid => buffer53_outs_valid,
      ins_ready => buffer53_outs_ready,
      clk => clk,
      rst => rst,
      outs => trunci4_outs,
      outs_valid => trunci4_outs_valid,
      outs_ready => trunci4_outs_ready
    );

  shli5 : entity work.shli(arch) generic map(32)
    port map(
      lhs => buffer41_outs,
      lhs_valid => buffer41_outs_valid,
      lhs_ready => buffer41_outs_ready,
      rhs => fork21_outs_1,
      rhs_valid => fork21_outs_1_valid,
      rhs_ready => fork21_outs_1_ready,
      clk => clk,
      rst => rst,
      result => shli5_result,
      result_valid => shli5_result_valid,
      result_ready => shli5_result_ready
    );

  buffer41 : entity work.tfifo(arch) generic map(1, 32)
    port map(
      ins => fork12_outs_1,
      ins_valid => fork12_outs_1_valid,
      ins_ready => fork12_outs_1_ready,
      clk => clk,
      rst => rst,
      outs => buffer41_outs,
      outs_valid => buffer41_outs_valid,
      outs_ready => buffer41_outs_ready
    );

  buffer54 : entity work.oehb(arch) generic map(32)
    port map(
      ins => shli5_result,
      ins_valid => shli5_result_valid,
      ins_ready => shli5_result_ready,
      clk => clk,
      rst => rst,
      outs => buffer54_outs,
      outs_valid => buffer54_outs_valid,
      outs_ready => buffer54_outs_ready
    );

  trunci5 : entity work.trunci(arch) generic map(32, 7)
    port map(
      ins => buffer54_outs,
      ins_valid => buffer54_outs_valid,
      ins_ready => buffer54_outs_ready,
      clk => clk,
      rst => rst,
      outs => trunci5_outs,
      outs_valid => trunci5_outs_valid,
      outs_ready => trunci5_outs_ready
    );

  addi29 : entity work.addi(arch) generic map(7)
    port map(
      lhs => trunci4_outs,
      lhs_valid => trunci4_outs_valid,
      lhs_ready => trunci4_outs_ready,
      rhs => trunci5_outs,
      rhs_valid => trunci5_outs_valid,
      rhs_ready => trunci5_outs_ready,
      clk => clk,
      rst => rst,
      result => addi29_result,
      result_valid => addi29_result_valid,
      result_ready => addi29_result_ready
    );

  buffer56 : entity work.oehb(arch) generic map(7)
    port map(
      ins => addi29_result,
      ins_valid => addi29_result_valid,
      ins_ready => addi29_result_ready,
      clk => clk,
      rst => rst,
      outs => buffer56_outs,
      outs_valid => buffer56_outs_valid,
      outs_ready => buffer56_outs_ready
    );

  addi5 : entity work.addi(arch) generic map(7)
    port map(
      lhs => extsi60_outs,
      lhs_valid => extsi60_outs_valid,
      lhs_ready => extsi60_outs_ready,
      rhs => buffer56_outs,
      rhs_valid => buffer56_outs_valid,
      rhs_ready => buffer56_outs_ready,
      clk => clk,
      rst => rst,
      result => addi5_result,
      result_valid => addi5_result_valid,
      result_ready => addi5_result_ready
    );

  load1 : entity work.load(arch) generic map(32, 7)
    port map(
      addrIn => addi5_result,
      addrIn_valid => addi5_result_valid,
      addrIn_ready => addi5_result_ready,
      dataFromMem => mem_controller9_ldData_0,
      dataFromMem_valid => mem_controller9_ldData_0_valid,
      dataFromMem_ready => mem_controller9_ldData_0_ready,
      clk => clk,
      rst => rst,
      addrOut => load1_addrOut,
      addrOut_valid => load1_addrOut_valid,
      addrOut_ready => load1_addrOut_ready,
      dataOut => load1_dataOut,
      dataOut_valid => load1_dataOut_valid,
      dataOut_ready => load1_dataOut_ready
    );

  muli0 : entity work.muli(arch) generic map(32)
    port map(
      lhs => load0_dataOut,
      lhs_valid => load0_dataOut_valid,
      lhs_ready => load0_dataOut_ready,
      rhs => load1_dataOut,
      rhs_valid => load1_dataOut_valid,
      rhs_ready => load1_dataOut_ready,
      clk => clk,
      rst => rst,
      result => muli0_result,
      result_valid => muli0_result_valid,
      result_ready => muli0_result_ready
    );

  shli6 : entity work.shli(arch) generic map(32)
    port map(
      lhs => buffer43_outs,
      lhs_valid => buffer43_outs_valid,
      lhs_ready => buffer43_outs_ready,
      rhs => buffer42_outs,
      rhs_valid => buffer42_outs_valid,
      rhs_ready => buffer42_outs_ready,
      clk => clk,
      rst => rst,
      result => shli6_result,
      result_valid => shli6_result_valid,
      result_ready => shli6_result_ready
    );

  buffer42 : entity work.tfifo(arch) generic map(3, 32)
    port map(
      ins => fork20_outs_2,
      ins_valid => fork20_outs_2_valid,
      ins_ready => fork20_outs_2_ready,
      clk => clk,
      rst => rst,
      outs => buffer42_outs,
      outs_valid => buffer42_outs_valid,
      outs_ready => buffer42_outs_ready
    );

  buffer43 : entity work.tfifo(arch) generic map(3, 32)
    port map(
      ins => fork14_outs_2,
      ins_valid => fork14_outs_2_valid,
      ins_ready => fork14_outs_2_ready,
      clk => clk,
      rst => rst,
      outs => buffer43_outs,
      outs_valid => buffer43_outs_valid,
      outs_ready => buffer43_outs_ready
    );

  shli7 : entity work.shli(arch) generic map(32)
    port map(
      lhs => buffer45_outs,
      lhs_valid => buffer45_outs_valid,
      lhs_ready => buffer45_outs_ready,
      rhs => buffer44_outs,
      rhs_valid => buffer44_outs_valid,
      rhs_ready => buffer44_outs_ready,
      clk => clk,
      rst => rst,
      result => shli7_result,
      result_valid => shli7_result_valid,
      result_ready => shli7_result_ready
    );

  buffer44 : entity work.tfifo(arch) generic map(3, 32)
    port map(
      ins => fork21_outs_2,
      ins_valid => fork21_outs_2_valid,
      ins_ready => fork21_outs_2_ready,
      clk => clk,
      rst => rst,
      outs => buffer44_outs,
      outs_valid => buffer44_outs_valid,
      outs_ready => buffer44_outs_ready
    );

  buffer45 : entity work.tfifo(arch) generic map(3, 32)
    port map(
      ins => fork14_outs_3,
      ins_valid => fork14_outs_3_valid,
      ins_ready => fork14_outs_3_ready,
      clk => clk,
      rst => rst,
      outs => buffer45_outs,
      outs_valid => buffer45_outs_valid,
      outs_ready => buffer45_outs_ready
    );

  buffer57 : entity work.oehb(arch) generic map(32)
    port map(
      ins => shli6_result,
      ins_valid => shli6_result_valid,
      ins_ready => shli6_result_ready,
      clk => clk,
      rst => rst,
      outs => buffer57_outs,
      outs_valid => buffer57_outs_valid,
      outs_ready => buffer57_outs_ready
    );

  buffer58 : entity work.oehb(arch) generic map(32)
    port map(
      ins => shli7_result,
      ins_valid => shli7_result_valid,
      ins_ready => shli7_result_ready,
      clk => clk,
      rst => rst,
      outs => buffer58_outs,
      outs_valid => buffer58_outs_valid,
      outs_ready => buffer58_outs_ready
    );

  addi30 : entity work.addi(arch) generic map(32)
    port map(
      lhs => buffer57_outs,
      lhs_valid => buffer57_outs_valid,
      lhs_ready => buffer57_outs_ready,
      rhs => buffer58_outs,
      rhs_valid => buffer58_outs_valid,
      rhs_ready => buffer58_outs_ready,
      clk => clk,
      rst => rst,
      result => addi30_result,
      result_valid => addi30_result_valid,
      result_ready => addi30_result_ready
    );

  buffer61 : entity work.oehb(arch) generic map(32)
    port map(
      ins => addi30_result,
      ins_valid => addi30_result_valid,
      ins_ready => addi30_result_ready,
      clk => clk,
      rst => rst,
      outs => buffer61_outs,
      outs_valid => buffer61_outs_valid,
      outs_ready => buffer61_outs_ready
    );

  addi6 : entity work.addi(arch) generic map(32)
    port map(
      lhs => buffer46_outs,
      lhs_valid => buffer46_outs_valid,
      lhs_ready => buffer46_outs_ready,
      rhs => buffer61_outs,
      rhs_valid => buffer61_outs_valid,
      rhs_ready => buffer61_outs_ready,
      clk => clk,
      rst => rst,
      result => addi6_result,
      result_valid => addi6_result_valid,
      result_ready => addi6_result_ready
    );

  buffer46 : entity work.tfifo(arch) generic map(3, 32)
    port map(
      ins => fork16_outs_0,
      ins_valid => fork16_outs_0_valid,
      ins_ready => fork16_outs_0_ready,
      clk => clk,
      rst => rst,
      outs => buffer46_outs,
      outs_valid => buffer46_outs_valid,
      outs_ready => buffer46_outs_ready
    );

  buffer25 : entity work.tehb_dataless(arch)
    port map(
      ins_valid => mux31_outs_valid,
      ins_ready => mux31_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer25_outs_valid,
      outs_ready => buffer25_outs_ready
    );

  gate0 : entity work.gate(arch) generic map(3, 32)
    port map(
      ins(0) => addi6_result,
      ins_valid(0) => addi6_result_valid,
      ins_valid(1) => fork10_outs_1_valid,
      ins_valid(2) => buffer25_outs_valid,
      ins_ready(0) => addi6_result_ready,
      ins_ready(1) => fork10_outs_1_ready,
      ins_ready(2) => buffer25_outs_ready,
      clk => clk,
      rst => rst,
      outs => gate0_outs,
      outs_valid => gate0_outs_valid,
      outs_ready => gate0_outs_ready
    );

  trunci6 : entity work.trunci(arch) generic map(32, 7)
    port map(
      ins => gate0_outs,
      ins_valid => gate0_outs_valid,
      ins_ready => gate0_outs_ready,
      clk => clk,
      rst => rst,
      outs => trunci6_outs,
      outs_valid => trunci6_outs_valid,
      outs_ready => trunci6_outs_ready
    );

  load2 : entity work.load(arch) generic map(32, 7)
    port map(
      addrIn => trunci6_outs,
      addrIn_valid => trunci6_outs_valid,
      addrIn_ready => trunci6_outs_ready,
      dataFromMem => mem_controller6_ldData_0,
      dataFromMem_valid => mem_controller6_ldData_0_valid,
      dataFromMem_ready => mem_controller6_ldData_0_ready,
      clk => clk,
      rst => rst,
      addrOut => load2_addrOut,
      addrOut_valid => load2_addrOut_valid,
      addrOut_ready => load2_addrOut_ready,
      dataOut => load2_dataOut,
      dataOut_valid => load2_dataOut_valid,
      dataOut_ready => load2_dataOut_ready
    );

  addi0 : entity work.addi(arch) generic map(32)
    port map(
      lhs => load2_dataOut,
      lhs_valid => load2_dataOut_valid,
      lhs_ready => load2_dataOut_ready,
      rhs => muli0_result,
      rhs_valid => muli0_result_valid,
      rhs_ready => muli0_result_ready,
      clk => clk,
      rst => rst,
      result => addi0_result,
      result_valid => addi0_result_valid,
      result_ready => addi0_result_ready
    );

  shli8 : entity work.shli(arch) generic map(32)
    port map(
      lhs => buffer48_outs,
      lhs_valid => buffer48_outs_valid,
      lhs_ready => buffer48_outs_ready,
      rhs => buffer47_outs,
      rhs_valid => buffer47_outs_valid,
      rhs_ready => buffer47_outs_ready,
      clk => clk,
      rst => rst,
      result => shli8_result,
      result_valid => shli8_result_valid,
      result_ready => shli8_result_ready
    );

  buffer47 : entity work.tfifo(arch) generic map(3, 32)
    port map(
      ins => fork20_outs_3,
      ins_valid => fork20_outs_3_valid,
      ins_ready => fork20_outs_3_ready,
      clk => clk,
      rst => rst,
      outs => buffer47_outs,
      outs_valid => buffer47_outs_valid,
      outs_ready => buffer47_outs_ready
    );

  buffer48 : entity work.tfifo(arch) generic map(3, 32)
    port map(
      ins => fork14_outs_4,
      ins_valid => fork14_outs_4_valid,
      ins_ready => fork14_outs_4_ready,
      clk => clk,
      rst => rst,
      outs => buffer48_outs,
      outs_valid => buffer48_outs_valid,
      outs_ready => buffer48_outs_ready
    );

  shli9 : entity work.shli(arch) generic map(32)
    port map(
      lhs => buffer50_outs,
      lhs_valid => buffer50_outs_valid,
      lhs_ready => buffer50_outs_ready,
      rhs => buffer49_outs,
      rhs_valid => buffer49_outs_valid,
      rhs_ready => buffer49_outs_ready,
      clk => clk,
      rst => rst,
      result => shli9_result,
      result_valid => shli9_result_valid,
      result_ready => shli9_result_ready
    );

  buffer49 : entity work.tfifo(arch) generic map(3, 32)
    port map(
      ins => fork21_outs_3,
      ins_valid => fork21_outs_3_valid,
      ins_ready => fork21_outs_3_ready,
      clk => clk,
      rst => rst,
      outs => buffer49_outs,
      outs_valid => buffer49_outs_valid,
      outs_ready => buffer49_outs_ready
    );

  buffer50 : entity work.tfifo(arch) generic map(3, 32)
    port map(
      ins => fork14_outs_5,
      ins_valid => fork14_outs_5_valid,
      ins_ready => fork14_outs_5_ready,
      clk => clk,
      rst => rst,
      outs => buffer50_outs,
      outs_valid => buffer50_outs_valid,
      outs_ready => buffer50_outs_ready
    );

  buffer62 : entity work.oehb(arch) generic map(32)
    port map(
      ins => shli8_result,
      ins_valid => shli8_result_valid,
      ins_ready => shli8_result_ready,
      clk => clk,
      rst => rst,
      outs => buffer62_outs,
      outs_valid => buffer62_outs_valid,
      outs_ready => buffer62_outs_ready
    );

  buffer63 : entity work.oehb(arch) generic map(32)
    port map(
      ins => shli9_result,
      ins_valid => shli9_result_valid,
      ins_ready => shli9_result_ready,
      clk => clk,
      rst => rst,
      outs => buffer63_outs,
      outs_valid => buffer63_outs_valid,
      outs_ready => buffer63_outs_ready
    );

  addi31 : entity work.addi(arch) generic map(32)
    port map(
      lhs => buffer62_outs,
      lhs_valid => buffer62_outs_valid,
      lhs_ready => buffer62_outs_ready,
      rhs => buffer63_outs,
      rhs_valid => buffer63_outs_valid,
      rhs_ready => buffer63_outs_ready,
      clk => clk,
      rst => rst,
      result => addi31_result,
      result_valid => addi31_result_valid,
      result_ready => addi31_result_ready
    );

  buffer64 : entity work.oehb(arch) generic map(32)
    port map(
      ins => addi31_result,
      ins_valid => addi31_result_valid,
      ins_ready => addi31_result_ready,
      clk => clk,
      rst => rst,
      outs => buffer64_outs,
      outs_valid => buffer64_outs_valid,
      outs_ready => buffer64_outs_ready
    );

  addi7 : entity work.addi(arch) generic map(32)
    port map(
      lhs => buffer51_outs,
      lhs_valid => buffer51_outs_valid,
      lhs_ready => buffer51_outs_ready,
      rhs => buffer64_outs,
      rhs_valid => buffer64_outs_valid,
      rhs_ready => buffer64_outs_ready,
      clk => clk,
      rst => rst,
      result => addi7_result,
      result_valid => addi7_result_valid,
      result_ready => addi7_result_ready
    );

  buffer51 : entity work.tfifo(arch) generic map(4, 32)
    port map(
      ins => fork16_outs_1,
      ins_valid => fork16_outs_1_valid,
      ins_ready => fork16_outs_1_ready,
      clk => clk,
      rst => rst,
      outs => buffer51_outs,
      outs_valid => buffer51_outs_valid,
      outs_ready => buffer51_outs_ready
    );

  buffer1 : entity work.tfifo_dataless(arch) generic map(1)
    port map(
      ins_valid => store1_doneOut_valid,
      ins_ready => store1_doneOut_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer1_outs_valid,
      outs_ready => buffer1_outs_ready
    );

  gate1 : entity work.gate(arch) generic map(2, 32)
    port map(
      ins(0) => addi7_result,
      ins_valid(0) => addi7_result_valid,
      ins_valid(1) => fork10_outs_0_valid,
      ins_ready(0) => addi7_result_ready,
      ins_ready(1) => fork10_outs_0_ready,
      clk => clk,
      rst => rst,
      outs => gate1_outs,
      outs_valid => gate1_outs_valid,
      outs_ready => gate1_outs_ready
    );

  trunci7 : entity work.trunci(arch) generic map(32, 7)
    port map(
      ins => gate1_outs,
      ins_valid => gate1_outs_valid,
      ins_ready => gate1_outs_ready,
      clk => clk,
      rst => rst,
      outs => trunci7_outs,
      outs_valid => trunci7_outs_valid,
      outs_ready => trunci7_outs_ready
    );

  store1 : entity work.store(arch) generic map(32, 7)
    port map(
      addrIn => trunci7_outs,
      addrIn_valid => trunci7_outs_valid,
      addrIn_ready => trunci7_outs_ready,
      dataIn => addi0_result,
      dataIn_valid => addi0_result_valid,
      dataIn_ready => addi0_result_ready,
      doneFromMem_valid => mem_controller6_stDone_1_valid,
      doneFromMem_ready => mem_controller6_stDone_1_ready,
      clk => clk,
      rst => rst,
      addrOut => store1_addrOut,
      addrOut_valid => store1_addrOut_valid,
      addrOut_ready => store1_addrOut_ready,
      dataToMem => store1_dataToMem,
      dataToMem_valid => store1_dataToMem_valid,
      dataToMem_ready => store1_dataToMem_ready,
      doneOut_valid => store1_doneOut_valid,
      doneOut_ready => store1_doneOut_ready
    );

  addi18 : entity work.addi(arch) generic map(6)
    port map(
      lhs => extsi57_outs,
      lhs_valid => extsi57_outs_valid,
      lhs_ready => extsi57_outs_ready,
      rhs => extsi63_outs,
      rhs_valid => extsi63_outs_valid,
      rhs_ready => extsi63_outs_ready,
      clk => clk,
      rst => rst,
      result => addi18_result,
      result_valid => addi18_result_valid,
      result_ready => addi18_result_ready
    );

  buffer67 : entity work.oehb(arch) generic map(6)
    port map(
      ins => addi18_result,
      ins_valid => addi18_result_valid,
      ins_ready => addi18_result_ready,
      clk => clk,
      rst => rst,
      outs => buffer67_outs,
      outs_valid => buffer67_outs_valid,
      outs_ready => buffer67_outs_ready
    );

  fork22 : entity work.handshake_fork(arch) generic map(2, 6)
    port map(
      ins => buffer67_outs,
      ins_valid => buffer67_outs_valid,
      ins_ready => buffer67_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork22_outs_0,
      outs(1) => fork22_outs_1,
      outs_valid(0) => fork22_outs_0_valid,
      outs_valid(1) => fork22_outs_1_valid,
      outs_ready(0) => fork22_outs_0_ready,
      outs_ready(1) => fork22_outs_1_ready
    );

  trunci8 : entity work.trunci(arch) generic map(6, 5)
    port map(
      ins => fork22_outs_0,
      ins_valid => fork22_outs_0_valid,
      ins_ready => fork22_outs_0_ready,
      clk => clk,
      rst => rst,
      outs => trunci8_outs,
      outs_valid => trunci8_outs_valid,
      outs_ready => trunci8_outs_ready
    );

  cmpi0 : entity work.handshake_cmpi_0(arch) generic map(6)
    port map(
      lhs => fork22_outs_1,
      lhs_valid => fork22_outs_1_valid,
      lhs_ready => fork22_outs_1_ready,
      rhs => extsi62_outs,
      rhs_valid => extsi62_outs_valid,
      rhs_ready => extsi62_outs_ready,
      clk => clk,
      rst => rst,
      result => cmpi0_result,
      result_valid => cmpi0_result_valid,
      result_ready => cmpi0_result_ready
    );

  buffer68 : entity work.oehb(arch) generic map(1)
    port map(
      ins => cmpi0_result,
      ins_valid => cmpi0_result_valid,
      ins_ready => cmpi0_result_ready,
      clk => clk,
      rst => rst,
      outs => buffer68_outs,
      outs_valid => buffer68_outs_valid,
      outs_ready => buffer68_outs_ready
    );

  fork23 : entity work.handshake_fork(arch) generic map(7, 1)
    port map(
      ins => buffer68_outs,
      ins_valid => buffer68_outs_valid,
      ins_ready => buffer68_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork23_outs_0,
      outs(1) => fork23_outs_1,
      outs(2) => fork23_outs_2,
      outs(3) => fork23_outs_3,
      outs(4) => fork23_outs_4,
      outs(5) => fork23_outs_5,
      outs(6) => fork23_outs_6,
      outs_valid(0) => fork23_outs_0_valid,
      outs_valid(1) => fork23_outs_1_valid,
      outs_valid(2) => fork23_outs_2_valid,
      outs_valid(3) => fork23_outs_3_valid,
      outs_valid(4) => fork23_outs_4_valid,
      outs_valid(5) => fork23_outs_5_valid,
      outs_valid(6) => fork23_outs_6_valid,
      outs_ready(0) => fork23_outs_0_ready,
      outs_ready(1) => fork23_outs_1_ready,
      outs_ready(2) => fork23_outs_2_ready,
      outs_ready(3) => fork23_outs_3_ready,
      outs_ready(4) => fork23_outs_4_ready,
      outs_ready(5) => fork23_outs_5_ready,
      outs_ready(6) => fork23_outs_6_ready
    );

  cond_br9 : entity work.cond_br(arch) generic map(5)
    port map(
      condition => fork23_outs_0,
      condition_valid => fork23_outs_0_valid,
      condition_ready => fork23_outs_0_ready,
      data => trunci8_outs,
      data_valid => trunci8_outs_valid,
      data_ready => trunci8_outs_ready,
      clk => clk,
      rst => rst,
      trueOut => cond_br9_trueOut,
      trueOut_valid => cond_br9_trueOut_valid,
      trueOut_ready => cond_br9_trueOut_ready,
      falseOut => cond_br9_falseOut,
      falseOut_valid => cond_br9_falseOut_valid,
      falseOut_ready => cond_br9_falseOut_ready
    );

  sink1 : entity work.sink(arch) generic map(5)
    port map(
      ins => cond_br9_falseOut,
      ins_valid => cond_br9_falseOut_valid,
      ins_ready => cond_br9_falseOut_ready,
      clk => clk,
      rst => rst
    );

  cond_br10 : entity work.cond_br(arch) generic map(5)
    port map(
      condition => buffer55_outs,
      condition_valid => buffer55_outs_valid,
      condition_ready => buffer55_outs_ready,
      data => fork13_outs_0,
      data_valid => fork13_outs_0_valid,
      data_ready => fork13_outs_0_ready,
      clk => clk,
      rst => rst,
      trueOut => cond_br10_trueOut,
      trueOut_valid => cond_br10_trueOut_valid,
      trueOut_ready => cond_br10_trueOut_ready,
      falseOut => cond_br10_falseOut,
      falseOut_valid => cond_br10_falseOut_valid,
      falseOut_ready => cond_br10_falseOut_ready
    );

  buffer55 : entity work.tfifo(arch) generic map(1, 1)
    port map(
      ins => fork23_outs_1,
      ins_valid => fork23_outs_1_valid,
      ins_ready => fork23_outs_1_ready,
      clk => clk,
      rst => rst,
      outs => buffer55_outs,
      outs_valid => buffer55_outs_valid,
      outs_ready => buffer55_outs_ready
    );

  cond_br11 : entity work.cond_br(arch) generic map(5)
    port map(
      condition => fork23_outs_2,
      condition_valid => fork23_outs_2_valid,
      condition_ready => fork23_outs_2_ready,
      data => fork15_outs_1,
      data_valid => fork15_outs_1_valid,
      data_ready => fork15_outs_1_ready,
      clk => clk,
      rst => rst,
      trueOut => cond_br11_trueOut,
      trueOut_valid => cond_br11_trueOut_valid,
      trueOut_ready => cond_br11_trueOut_ready,
      falseOut => cond_br11_falseOut,
      falseOut_valid => cond_br11_falseOut_valid,
      falseOut_ready => cond_br11_falseOut_ready
    );

  buffer36 : entity work.oehb_dataless(arch)
    port map(
      ins_valid => fork18_outs_1_valid,
      ins_ready => fork18_outs_1_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer36_outs_valid,
      outs_ready => buffer36_outs_ready
    );

  cond_br12 : entity work.cond_br_dataless(arch)
    port map(
      condition => buffer59_outs,
      condition_valid => buffer59_outs_valid,
      condition_ready => buffer59_outs_ready,
      data_valid => buffer36_outs_valid,
      data_ready => buffer36_outs_ready,
      clk => clk,
      rst => rst,
      trueOut_valid => cond_br12_trueOut_valid,
      trueOut_ready => cond_br12_trueOut_ready,
      falseOut_valid => cond_br12_falseOut_valid,
      falseOut_ready => cond_br12_falseOut_ready
    );

  buffer59 : entity work.tfifo(arch) generic map(1, 1)
    port map(
      ins => fork23_outs_6,
      ins_valid => fork23_outs_6_valid,
      ins_ready => fork23_outs_6_ready,
      clk => clk,
      rst => rst,
      outs => buffer59_outs,
      outs_valid => buffer59_outs_valid,
      outs_ready => buffer59_outs_ready
    );

  cond_br118 : entity work.cond_br_dataless(arch)
    port map(
      condition => buffer60_outs,
      condition_valid => buffer60_outs_valid,
      condition_ready => buffer60_outs_ready,
      data_valid => cond_br116_falseOut_valid,
      data_ready => cond_br116_falseOut_ready,
      clk => clk,
      rst => rst,
      trueOut_valid => cond_br118_trueOut_valid,
      trueOut_ready => cond_br118_trueOut_ready,
      falseOut_valid => cond_br118_falseOut_valid,
      falseOut_ready => cond_br118_falseOut_ready
    );

  buffer60 : entity work.tfifo(arch) generic map(1, 1)
    port map(
      ins => fork25_outs_3,
      ins_valid => fork25_outs_3_valid,
      ins_ready => fork25_outs_3_ready,
      clk => clk,
      rst => rst,
      outs => buffer60_outs,
      outs_valid => buffer60_outs_valid,
      outs_ready => buffer60_outs_ready
    );

  cond_br119 : entity work.cond_br_dataless(arch)
    port map(
      condition => fork25_outs_2,
      condition_valid => fork25_outs_2_valid,
      condition_ready => fork25_outs_2_ready,
      data_valid => fork8_outs_0_valid,
      data_ready => fork8_outs_0_ready,
      clk => clk,
      rst => rst,
      trueOut_valid => cond_br119_trueOut_valid,
      trueOut_ready => cond_br119_trueOut_ready,
      falseOut_valid => cond_br119_falseOut_valid,
      falseOut_ready => cond_br119_falseOut_ready
    );

  sink2 : entity work.sink_dataless(arch)
    port map(
      ins_valid => cond_br119_trueOut_valid,
      ins_ready => cond_br119_trueOut_ready,
      clk => clk,
      rst => rst
    );

  extsi64 : entity work.extsi(arch) generic map(5, 6)
    port map(
      ins => cond_br11_falseOut,
      ins_valid => cond_br11_falseOut_valid,
      ins_ready => cond_br11_falseOut_ready,
      clk => clk,
      rst => rst,
      outs => extsi64_outs,
      outs_valid => extsi64_outs_valid,
      outs_ready => extsi64_outs_ready
    );

  source5 : entity work.source(arch)
    port map(
      clk => clk,
      rst => rst,
      outs_valid => source5_outs_valid,
      outs_ready => source5_outs_ready
    );

  constant55 : entity work.handshake_constant_3(arch) generic map(5)
    port map(
      ctrl_valid => source5_outs_valid,
      ctrl_ready => source5_outs_ready,
      clk => clk,
      rst => rst,
      outs => constant55_outs,
      outs_valid => constant55_outs_valid,
      outs_ready => constant55_outs_ready
    );

  extsi65 : entity work.extsi(arch) generic map(5, 6)
    port map(
      ins => constant55_outs,
      ins_valid => constant55_outs_valid,
      ins_ready => constant55_outs_ready,
      clk => clk,
      rst => rst,
      outs => extsi65_outs,
      outs_valid => extsi65_outs_valid,
      outs_ready => extsi65_outs_ready
    );

  source6 : entity work.source(arch)
    port map(
      clk => clk,
      rst => rst,
      outs_valid => source6_outs_valid,
      outs_ready => source6_outs_ready
    );

  constant56 : entity work.handshake_constant_1(arch) generic map(2)
    port map(
      ctrl_valid => source6_outs_valid,
      ctrl_ready => source6_outs_ready,
      clk => clk,
      rst => rst,
      outs => constant56_outs,
      outs_valid => constant56_outs_valid,
      outs_ready => constant56_outs_ready
    );

  extsi66 : entity work.extsi(arch) generic map(2, 6)
    port map(
      ins => constant56_outs,
      ins_valid => constant56_outs_valid,
      ins_ready => constant56_outs_ready,
      clk => clk,
      rst => rst,
      outs => extsi66_outs,
      outs_valid => extsi66_outs_valid,
      outs_ready => extsi66_outs_ready
    );

  addi19 : entity work.addi(arch) generic map(6)
    port map(
      lhs => extsi64_outs,
      lhs_valid => extsi64_outs_valid,
      lhs_ready => extsi64_outs_ready,
      rhs => extsi66_outs,
      rhs_valid => extsi66_outs_valid,
      rhs_ready => extsi66_outs_ready,
      clk => clk,
      rst => rst,
      result => addi19_result,
      result_valid => addi19_result_valid,
      result_ready => addi19_result_ready
    );

  buffer69 : entity work.oehb(arch) generic map(6)
    port map(
      ins => addi19_result,
      ins_valid => addi19_result_valid,
      ins_ready => addi19_result_ready,
      clk => clk,
      rst => rst,
      outs => buffer69_outs,
      outs_valid => buffer69_outs_valid,
      outs_ready => buffer69_outs_ready
    );

  fork24 : entity work.handshake_fork(arch) generic map(2, 6)
    port map(
      ins => buffer69_outs,
      ins_valid => buffer69_outs_valid,
      ins_ready => buffer69_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork24_outs_0,
      outs(1) => fork24_outs_1,
      outs_valid(0) => fork24_outs_0_valid,
      outs_valid(1) => fork24_outs_1_valid,
      outs_ready(0) => fork24_outs_0_ready,
      outs_ready(1) => fork24_outs_1_ready
    );

  trunci9 : entity work.trunci(arch) generic map(6, 5)
    port map(
      ins => fork24_outs_0,
      ins_valid => fork24_outs_0_valid,
      ins_ready => fork24_outs_0_ready,
      clk => clk,
      rst => rst,
      outs => trunci9_outs,
      outs_valid => trunci9_outs_valid,
      outs_ready => trunci9_outs_ready
    );

  cmpi1 : entity work.handshake_cmpi_0(arch) generic map(6)
    port map(
      lhs => fork24_outs_1,
      lhs_valid => fork24_outs_1_valid,
      lhs_ready => fork24_outs_1_ready,
      rhs => extsi65_outs,
      rhs_valid => extsi65_outs_valid,
      rhs_ready => extsi65_outs_ready,
      clk => clk,
      rst => rst,
      result => cmpi1_result,
      result_valid => cmpi1_result_valid,
      result_ready => cmpi1_result_ready
    );

  buffer70 : entity work.oehb(arch) generic map(1)
    port map(
      ins => cmpi1_result,
      ins_valid => cmpi1_result_valid,
      ins_ready => cmpi1_result_ready,
      clk => clk,
      rst => rst,
      outs => buffer70_outs,
      outs_valid => buffer70_outs_valid,
      outs_ready => buffer70_outs_ready
    );

  fork25 : entity work.handshake_fork(arch) generic map(6, 1)
    port map(
      ins => buffer70_outs,
      ins_valid => buffer70_outs_valid,
      ins_ready => buffer70_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork25_outs_0,
      outs(1) => fork25_outs_1,
      outs(2) => fork25_outs_2,
      outs(3) => fork25_outs_3,
      outs(4) => fork25_outs_4,
      outs(5) => fork25_outs_5,
      outs_valid(0) => fork25_outs_0_valid,
      outs_valid(1) => fork25_outs_1_valid,
      outs_valid(2) => fork25_outs_2_valid,
      outs_valid(3) => fork25_outs_3_valid,
      outs_valid(4) => fork25_outs_4_valid,
      outs_valid(5) => fork25_outs_5_valid,
      outs_ready(0) => fork25_outs_0_ready,
      outs_ready(1) => fork25_outs_1_ready,
      outs_ready(2) => fork25_outs_2_ready,
      outs_ready(3) => fork25_outs_3_ready,
      outs_ready(4) => fork25_outs_4_ready,
      outs_ready(5) => fork25_outs_5_ready
    );

  cond_br13 : entity work.cond_br(arch) generic map(5)
    port map(
      condition => fork25_outs_0,
      condition_valid => fork25_outs_0_valid,
      condition_ready => fork25_outs_0_ready,
      data => trunci9_outs,
      data_valid => trunci9_outs_valid,
      data_ready => trunci9_outs_ready,
      clk => clk,
      rst => rst,
      trueOut => cond_br13_trueOut,
      trueOut_valid => cond_br13_trueOut_valid,
      trueOut_ready => cond_br13_trueOut_ready,
      falseOut => cond_br13_falseOut,
      falseOut_valid => cond_br13_falseOut_valid,
      falseOut_ready => cond_br13_falseOut_ready
    );

  sink4 : entity work.sink(arch) generic map(5)
    port map(
      ins => cond_br13_falseOut,
      ins_valid => cond_br13_falseOut_valid,
      ins_ready => cond_br13_falseOut_ready,
      clk => clk,
      rst => rst
    );

  cond_br14 : entity work.cond_br(arch) generic map(5)
    port map(
      condition => fork25_outs_1,
      condition_valid => fork25_outs_1_valid,
      condition_ready => fork25_outs_1_ready,
      data => cond_br10_falseOut,
      data_valid => cond_br10_falseOut_valid,
      data_ready => cond_br10_falseOut_ready,
      clk => clk,
      rst => rst,
      trueOut => cond_br14_trueOut,
      trueOut_valid => cond_br14_trueOut_valid,
      trueOut_ready => cond_br14_trueOut_ready,
      falseOut => cond_br14_falseOut,
      falseOut_valid => cond_br14_falseOut_valid,
      falseOut_ready => cond_br14_falseOut_ready
    );

  cond_br15 : entity work.cond_br_dataless(arch)
    port map(
      condition => buffer66_outs,
      condition_valid => buffer66_outs_valid,
      condition_ready => buffer66_outs_ready,
      data_valid => cond_br12_falseOut_valid,
      data_ready => cond_br12_falseOut_ready,
      clk => clk,
      rst => rst,
      trueOut_valid => cond_br15_trueOut_valid,
      trueOut_ready => cond_br15_trueOut_ready,
      falseOut_valid => cond_br15_falseOut_valid,
      falseOut_ready => cond_br15_falseOut_ready
    );

  buffer66 : entity work.tfifo(arch) generic map(1, 1)
    port map(
      ins => fork25_outs_5,
      ins_valid => fork25_outs_5_valid,
      ins_ready => fork25_outs_5_ready,
      clk => clk,
      rst => rst,
      outs => buffer66_outs,
      outs_valid => buffer66_outs_valid,
      outs_ready => buffer66_outs_ready
    );

  cond_br120 : entity work.cond_br_dataless(arch)
    port map(
      condition => fork28_outs_2,
      condition_valid => fork28_outs_2_valid,
      condition_ready => fork28_outs_2_ready,
      data_valid => cond_br118_falseOut_valid,
      data_ready => cond_br118_falseOut_ready,
      clk => clk,
      rst => rst,
      trueOut_valid => cond_br120_trueOut_valid,
      trueOut_ready => cond_br120_trueOut_ready,
      falseOut_valid => cond_br120_falseOut_valid,
      falseOut_ready => cond_br120_falseOut_ready
    );

  cond_br121 : entity work.cond_br_dataless(arch)
    port map(
      condition => fork28_outs_1,
      condition_valid => fork28_outs_1_valid,
      condition_ready => fork28_outs_1_ready,
      data_valid => cond_br119_falseOut_valid,
      data_ready => cond_br119_falseOut_ready,
      clk => clk,
      rst => rst,
      trueOut_valid => cond_br121_trueOut_valid,
      trueOut_ready => cond_br121_trueOut_ready,
      falseOut_valid => cond_br121_falseOut_valid,
      falseOut_ready => cond_br121_falseOut_ready
    );

  sink5 : entity work.sink_dataless(arch)
    port map(
      ins_valid => cond_br121_trueOut_valid,
      ins_ready => cond_br121_trueOut_ready,
      clk => clk,
      rst => rst
    );

  buffer71 : entity work.oehb(arch) generic map(5)
    port map(
      ins => cond_br14_falseOut,
      ins_valid => cond_br14_falseOut_valid,
      ins_ready => cond_br14_falseOut_ready,
      clk => clk,
      rst => rst,
      outs => buffer71_outs,
      outs_valid => buffer71_outs_valid,
      outs_ready => buffer71_outs_ready
    );

  extsi67 : entity work.extsi(arch) generic map(5, 6)
    port map(
      ins => buffer71_outs,
      ins_valid => buffer71_outs_valid,
      ins_ready => buffer71_outs_ready,
      clk => clk,
      rst => rst,
      outs => extsi67_outs,
      outs_valid => extsi67_outs_valid,
      outs_ready => extsi67_outs_ready
    );

  fork26 : entity work.fork_dataless(arch) generic map(2)
    port map(
      ins_valid => cond_br15_falseOut_valid,
      ins_ready => cond_br15_falseOut_ready,
      clk => clk,
      rst => rst,
      outs_valid(0) => fork26_outs_0_valid,
      outs_valid(1) => fork26_outs_1_valid,
      outs_ready(0) => fork26_outs_0_ready,
      outs_ready(1) => fork26_outs_1_ready
    );

  constant57 : entity work.handshake_constant_0(arch) generic map(1)
    port map(
      ctrl_valid => fork26_outs_0_valid,
      ctrl_ready => fork26_outs_0_ready,
      clk => clk,
      rst => rst,
      outs => constant57_outs,
      outs_valid => constant57_outs_valid,
      outs_ready => constant57_outs_ready
    );

  source7 : entity work.source(arch)
    port map(
      clk => clk,
      rst => rst,
      outs_valid => source7_outs_valid,
      outs_ready => source7_outs_ready
    );

  constant58 : entity work.handshake_constant_3(arch) generic map(5)
    port map(
      ctrl_valid => source7_outs_valid,
      ctrl_ready => source7_outs_ready,
      clk => clk,
      rst => rst,
      outs => constant58_outs,
      outs_valid => constant58_outs_valid,
      outs_ready => constant58_outs_ready
    );

  extsi68 : entity work.extsi(arch) generic map(5, 6)
    port map(
      ins => constant58_outs,
      ins_valid => constant58_outs_valid,
      ins_ready => constant58_outs_ready,
      clk => clk,
      rst => rst,
      outs => extsi68_outs,
      outs_valid => extsi68_outs_valid,
      outs_ready => extsi68_outs_ready
    );

  source8 : entity work.source(arch)
    port map(
      clk => clk,
      rst => rst,
      outs_valid => source8_outs_valid,
      outs_ready => source8_outs_ready
    );

  constant59 : entity work.handshake_constant_1(arch) generic map(2)
    port map(
      ctrl_valid => source8_outs_valid,
      ctrl_ready => source8_outs_ready,
      clk => clk,
      rst => rst,
      outs => constant59_outs,
      outs_valid => constant59_outs_valid,
      outs_ready => constant59_outs_ready
    );

  extsi69 : entity work.extsi(arch) generic map(2, 6)
    port map(
      ins => constant59_outs,
      ins_valid => constant59_outs_valid,
      ins_ready => constant59_outs_ready,
      clk => clk,
      rst => rst,
      outs => extsi69_outs,
      outs_valid => extsi69_outs_valid,
      outs_ready => extsi69_outs_ready
    );

  addi20 : entity work.addi(arch) generic map(6)
    port map(
      lhs => extsi67_outs,
      lhs_valid => extsi67_outs_valid,
      lhs_ready => extsi67_outs_ready,
      rhs => extsi69_outs,
      rhs_valid => extsi69_outs_valid,
      rhs_ready => extsi69_outs_ready,
      clk => clk,
      rst => rst,
      result => addi20_result,
      result_valid => addi20_result_valid,
      result_ready => addi20_result_ready
    );

  buffer72 : entity work.oehb(arch) generic map(6)
    port map(
      ins => addi20_result,
      ins_valid => addi20_result_valid,
      ins_ready => addi20_result_ready,
      clk => clk,
      rst => rst,
      outs => buffer72_outs,
      outs_valid => buffer72_outs_valid,
      outs_ready => buffer72_outs_ready
    );

  fork27 : entity work.handshake_fork(arch) generic map(2, 6)
    port map(
      ins => buffer72_outs,
      ins_valid => buffer72_outs_valid,
      ins_ready => buffer72_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork27_outs_0,
      outs(1) => fork27_outs_1,
      outs_valid(0) => fork27_outs_0_valid,
      outs_valid(1) => fork27_outs_1_valid,
      outs_ready(0) => fork27_outs_0_ready,
      outs_ready(1) => fork27_outs_1_ready
    );

  trunci10 : entity work.trunci(arch) generic map(6, 5)
    port map(
      ins => fork27_outs_0,
      ins_valid => fork27_outs_0_valid,
      ins_ready => fork27_outs_0_ready,
      clk => clk,
      rst => rst,
      outs => trunci10_outs,
      outs_valid => trunci10_outs_valid,
      outs_ready => trunci10_outs_ready
    );

  cmpi2 : entity work.handshake_cmpi_0(arch) generic map(6)
    port map(
      lhs => fork27_outs_1,
      lhs_valid => fork27_outs_1_valid,
      lhs_ready => fork27_outs_1_ready,
      rhs => extsi68_outs,
      rhs_valid => extsi68_outs_valid,
      rhs_ready => extsi68_outs_ready,
      clk => clk,
      rst => rst,
      result => cmpi2_result,
      result_valid => cmpi2_result_valid,
      result_ready => cmpi2_result_ready
    );

  buffer73 : entity work.oehb(arch) generic map(1)
    port map(
      ins => cmpi2_result,
      ins_valid => cmpi2_result_valid,
      ins_ready => cmpi2_result_ready,
      clk => clk,
      rst => rst,
      outs => buffer73_outs,
      outs_valid => buffer73_outs_valid,
      outs_ready => buffer73_outs_ready
    );

  fork28 : entity work.handshake_fork(arch) generic map(6, 1)
    port map(
      ins => buffer73_outs,
      ins_valid => buffer73_outs_valid,
      ins_ready => buffer73_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork28_outs_0,
      outs(1) => fork28_outs_1,
      outs(2) => fork28_outs_2,
      outs(3) => fork28_outs_3,
      outs(4) => fork28_outs_4,
      outs(5) => fork28_outs_5,
      outs_valid(0) => fork28_outs_0_valid,
      outs_valid(1) => fork28_outs_1_valid,
      outs_valid(2) => fork28_outs_2_valid,
      outs_valid(3) => fork28_outs_3_valid,
      outs_valid(4) => fork28_outs_4_valid,
      outs_valid(5) => fork28_outs_5_valid,
      outs_ready(0) => fork28_outs_0_ready,
      outs_ready(1) => fork28_outs_1_ready,
      outs_ready(2) => fork28_outs_2_ready,
      outs_ready(3) => fork28_outs_3_ready,
      outs_ready(4) => fork28_outs_4_ready,
      outs_ready(5) => fork28_outs_5_ready
    );

  cond_br16 : entity work.cond_br(arch) generic map(5)
    port map(
      condition => fork28_outs_0,
      condition_valid => fork28_outs_0_valid,
      condition_ready => fork28_outs_0_ready,
      data => trunci10_outs,
      data_valid => trunci10_outs_valid,
      data_ready => trunci10_outs_ready,
      clk => clk,
      rst => rst,
      trueOut => cond_br16_trueOut,
      trueOut_valid => cond_br16_trueOut_valid,
      trueOut_ready => cond_br16_trueOut_ready,
      falseOut => cond_br16_falseOut,
      falseOut_valid => cond_br16_falseOut_valid,
      falseOut_ready => cond_br16_falseOut_ready
    );

  sink7 : entity work.sink(arch) generic map(5)
    port map(
      ins => cond_br16_falseOut,
      ins_valid => cond_br16_falseOut_valid,
      ins_ready => cond_br16_falseOut_ready,
      clk => clk,
      rst => rst
    );

  cond_br17 : entity work.cond_br_dataless(arch)
    port map(
      condition => fork28_outs_4,
      condition_valid => fork28_outs_4_valid,
      condition_ready => fork28_outs_4_ready,
      data_valid => fork26_outs_1_valid,
      data_ready => fork26_outs_1_ready,
      clk => clk,
      rst => rst,
      trueOut_valid => cond_br17_trueOut_valid,
      trueOut_ready => cond_br17_trueOut_ready,
      falseOut_valid => cond_br17_falseOut_valid,
      falseOut_ready => cond_br17_falseOut_ready
    );

  cond_br18 : entity work.cond_br(arch) generic map(1)
    port map(
      condition => fork28_outs_5,
      condition_valid => fork28_outs_5_valid,
      condition_ready => fork28_outs_5_ready,
      data => constant57_outs,
      data_valid => constant57_outs_valid,
      data_ready => constant57_outs_ready,
      clk => clk,
      rst => rst,
      trueOut => cond_br18_trueOut,
      trueOut_valid => cond_br18_trueOut_valid,
      trueOut_ready => cond_br18_trueOut_ready,
      falseOut => cond_br18_falseOut,
      falseOut_valid => cond_br18_falseOut_valid,
      falseOut_ready => cond_br18_falseOut_ready
    );

  sink8 : entity work.sink(arch) generic map(1)
    port map(
      ins => cond_br18_trueOut,
      ins_valid => cond_br18_trueOut_valid,
      ins_ready => cond_br18_trueOut_ready,
      clk => clk,
      rst => rst
    );

  extsi50 : entity work.extsi(arch) generic map(1, 5)
    port map(
      ins => cond_br18_falseOut,
      ins_valid => cond_br18_falseOut_valid,
      ins_ready => cond_br18_falseOut_ready,
      clk => clk,
      rst => rst,
      outs => extsi50_outs,
      outs_valid => extsi50_outs_valid,
      outs_ready => extsi50_outs_ready
    );

  mux35 : entity work.mux_dataless(arch) generic map(2, 1)
    port map(
      index => init14_outs,
      index_valid => init14_outs_valid,
      index_ready => init14_outs_ready,
      ins_valid(0) => fork0_outs_3_valid,
      ins_valid(1) => cond_br127_trueOut_valid,
      ins_ready(0) => fork0_outs_3_ready,
      ins_ready(1) => cond_br127_trueOut_ready,
      clk => clk,
      rst => rst,
      outs_valid => mux35_outs_valid,
      outs_ready => mux35_outs_ready
    );

  init14 : entity work.tehb_init(arch) generic map(1, 0)
    port map(
      ins => fork56_outs_3,
      ins_valid => fork56_outs_3_valid,
      ins_ready => fork56_outs_3_ready,
      clk => clk,
      rst => rst,
      outs => init14_outs,
      outs_valid => init14_outs_valid,
      outs_ready => init14_outs_ready
    );

  mux6 : entity work.mux(arch) generic map(2, 5, 1)
    port map(
      index => control_merge5_index,
      index_valid => control_merge5_index_valid,
      index_ready => control_merge5_index_ready,
      ins(0) => extsi50_outs,
      ins(1) => cond_br26_trueOut,
      ins_valid(0) => extsi50_outs_valid,
      ins_valid(1) => cond_br26_trueOut_valid,
      ins_ready(0) => extsi50_outs_ready,
      ins_ready(1) => cond_br26_trueOut_ready,
      clk => clk,
      rst => rst,
      outs => mux6_outs,
      outs_valid => mux6_outs_valid,
      outs_ready => mux6_outs_ready
    );

  control_merge5 : entity work.control_merge_dataless(arch) generic map(2, 1)
    port map(
      ins_valid(0) => cond_br17_falseOut_valid,
      ins_valid(1) => cond_br27_trueOut_valid,
      ins_ready(0) => cond_br17_falseOut_ready,
      ins_ready(1) => cond_br27_trueOut_ready,
      clk => clk,
      rst => rst,
      outs_valid => control_merge5_outs_valid,
      outs_ready => control_merge5_outs_ready,
      index => control_merge5_index,
      index_valid => control_merge5_index_valid,
      index_ready => control_merge5_index_ready
    );

  fork29 : entity work.fork_dataless(arch) generic map(2)
    port map(
      ins_valid => control_merge5_outs_valid,
      ins_ready => control_merge5_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid(0) => fork29_outs_0_valid,
      outs_valid(1) => fork29_outs_1_valid,
      outs_ready(0) => fork29_outs_0_ready,
      outs_ready(1) => fork29_outs_1_ready
    );

  constant60 : entity work.handshake_constant_0(arch) generic map(1)
    port map(
      ctrl_valid => fork29_outs_0_valid,
      ctrl_ready => fork29_outs_0_ready,
      clk => clk,
      rst => rst,
      outs => constant60_outs,
      outs_valid => constant60_outs_valid,
      outs_ready => constant60_outs_ready
    );

  extsi49 : entity work.extsi(arch) generic map(1, 5)
    port map(
      ins => constant60_outs,
      ins_valid => constant60_outs_valid,
      ins_ready => constant60_outs_ready,
      clk => clk,
      rst => rst,
      outs => extsi49_outs,
      outs_valid => extsi49_outs_valid,
      outs_ready => extsi49_outs_ready
    );

  buffer75 : entity work.tehb(arch) generic map(5)
    port map(
      ins => mux6_outs,
      ins_valid => mux6_outs_valid,
      ins_ready => mux6_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer75_outs,
      outs_valid => buffer75_outs_valid,
      outs_ready => buffer75_outs_ready
    );

  buffer74 : entity work.tehb_dataless(arch)
    port map(
      ins_valid => mux35_outs_valid,
      ins_ready => mux35_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer74_outs_valid,
      outs_ready => buffer74_outs_ready
    );

  mux40 : entity work.mux_dataless(arch) generic map(2, 1)
    port map(
      index => init19_outs,
      index_valid => init19_outs_valid,
      index_ready => init19_outs_ready,
      ins_valid(0) => buffer74_outs_valid,
      ins_valid(1) => cond_br125_trueOut_valid,
      ins_ready(0) => buffer74_outs_ready,
      ins_ready(1) => cond_br125_trueOut_ready,
      clk => clk,
      rst => rst,
      outs_valid => mux40_outs_valid,
      outs_ready => mux40_outs_ready
    );

  init19 : entity work.tehb_init(arch) generic map(1, 0)
    port map(
      ins => fork53_outs_4,
      ins_valid => fork53_outs_4_valid,
      ins_ready => fork53_outs_4_ready,
      clk => clk,
      rst => rst,
      outs => init19_outs,
      outs_valid => init19_outs_valid,
      outs_ready => init19_outs_ready
    );

  mux7 : entity work.mux(arch) generic map(2, 5, 1)
    port map(
      index => fork33_outs_1,
      index_valid => fork33_outs_1_valid,
      index_ready => fork33_outs_1_ready,
      ins(0) => extsi49_outs,
      ins(1) => cond_br23_trueOut,
      ins_valid(0) => extsi49_outs_valid,
      ins_valid(1) => cond_br23_trueOut_valid,
      ins_ready(0) => extsi49_outs_ready,
      ins_ready(1) => cond_br23_trueOut_ready,
      clk => clk,
      rst => rst,
      outs => mux7_outs,
      outs_valid => mux7_outs_valid,
      outs_ready => mux7_outs_ready
    );

  buffer78 : entity work.tehb(arch) generic map(5)
    port map(
      ins => mux7_outs,
      ins_valid => mux7_outs_valid,
      ins_ready => mux7_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer78_outs,
      outs_valid => buffer78_outs_valid,
      outs_ready => buffer78_outs_ready
    );

  fork30 : entity work.handshake_fork(arch) generic map(2, 5)
    port map(
      ins => buffer78_outs,
      ins_valid => buffer78_outs_valid,
      ins_ready => buffer78_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork30_outs_0,
      outs(1) => fork30_outs_1,
      outs_valid(0) => fork30_outs_0_valid,
      outs_valid(1) => fork30_outs_1_valid,
      outs_ready(0) => fork30_outs_0_ready,
      outs_ready(1) => fork30_outs_1_ready
    );

  extsi70 : entity work.extsi(arch) generic map(5, 7)
    port map(
      ins => fork30_outs_0,
      ins_valid => fork30_outs_0_valid,
      ins_ready => fork30_outs_0_ready,
      clk => clk,
      rst => rst,
      outs => extsi70_outs,
      outs_valid => extsi70_outs_valid,
      outs_ready => extsi70_outs_ready
    );

  mux8 : entity work.mux(arch) generic map(2, 5, 1)
    port map(
      index => fork33_outs_0,
      index_valid => fork33_outs_0_valid,
      index_ready => fork33_outs_0_ready,
      ins(0) => buffer75_outs,
      ins(1) => cond_br24_trueOut,
      ins_valid(0) => buffer75_outs_valid,
      ins_valid(1) => cond_br24_trueOut_valid,
      ins_ready(0) => buffer75_outs_ready,
      ins_ready(1) => cond_br24_trueOut_ready,
      clk => clk,
      rst => rst,
      outs => mux8_outs,
      outs_valid => mux8_outs_valid,
      outs_ready => mux8_outs_ready
    );

  buffer79 : entity work.oehb(arch) generic map(5)
    port map(
      ins => mux8_outs,
      ins_valid => mux8_outs_valid,
      ins_ready => mux8_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer79_outs,
      outs_valid => buffer79_outs_valid,
      outs_ready => buffer79_outs_ready
    );

  buffer80 : entity work.tehb(arch) generic map(5)
    port map(
      ins => buffer79_outs,
      ins_valid => buffer79_outs_valid,
      ins_ready => buffer79_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer80_outs,
      outs_valid => buffer80_outs_valid,
      outs_ready => buffer80_outs_ready
    );

  fork31 : entity work.handshake_fork(arch) generic map(2, 5)
    port map(
      ins => buffer80_outs,
      ins_valid => buffer80_outs_valid,
      ins_ready => buffer80_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork31_outs_0,
      outs(1) => fork31_outs_1,
      outs_valid(0) => fork31_outs_0_valid,
      outs_valid(1) => fork31_outs_1_valid,
      outs_ready(0) => fork31_outs_0_ready,
      outs_ready(1) => fork31_outs_1_ready
    );

  extsi71 : entity work.extsi(arch) generic map(5, 32)
    port map(
      ins => fork31_outs_1,
      ins_valid => fork31_outs_1_valid,
      ins_ready => fork31_outs_1_ready,
      clk => clk,
      rst => rst,
      outs => extsi71_outs,
      outs_valid => extsi71_outs_valid,
      outs_ready => extsi71_outs_ready
    );

  fork32 : entity work.handshake_fork(arch) generic map(2, 32)
    port map(
      ins => extsi71_outs,
      ins_valid => extsi71_outs_valid,
      ins_ready => extsi71_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork32_outs_0,
      outs(1) => fork32_outs_1,
      outs_valid(0) => fork32_outs_0_valid,
      outs_valid(1) => fork32_outs_1_valid,
      outs_ready(0) => fork32_outs_0_ready,
      outs_ready(1) => fork32_outs_1_ready
    );

  control_merge6 : entity work.control_merge_dataless(arch) generic map(2, 1)
    port map(
      ins_valid(0) => fork29_outs_1_valid,
      ins_valid(1) => cond_br25_trueOut_valid,
      ins_ready(0) => fork29_outs_1_ready,
      ins_ready(1) => cond_br25_trueOut_ready,
      clk => clk,
      rst => rst,
      outs_valid => control_merge6_outs_valid,
      outs_ready => control_merge6_outs_ready,
      index => control_merge6_index,
      index_valid => control_merge6_index_valid,
      index_ready => control_merge6_index_ready
    );

  fork33 : entity work.handshake_fork(arch) generic map(2, 1)
    port map(
      ins => control_merge6_index,
      ins_valid => control_merge6_index_valid,
      ins_ready => control_merge6_index_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork33_outs_0,
      outs(1) => fork33_outs_1,
      outs_valid(0) => fork33_outs_0_valid,
      outs_valid(1) => fork33_outs_1_valid,
      outs_ready(0) => fork33_outs_0_ready,
      outs_ready(1) => fork33_outs_1_ready
    );

  fork34 : entity work.fork_dataless(arch) generic map(3)
    port map(
      ins_valid => control_merge6_outs_valid,
      ins_ready => control_merge6_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid(0) => fork34_outs_0_valid,
      outs_valid(1) => fork34_outs_1_valid,
      outs_valid(2) => fork34_outs_2_valid,
      outs_ready(0) => fork34_outs_0_ready,
      outs_ready(1) => fork34_outs_1_ready,
      outs_ready(2) => fork34_outs_2_ready
    );

  constant61 : entity work.handshake_constant_1(arch) generic map(2)
    port map(
      ctrl_valid => fork34_outs_1_valid,
      ctrl_ready => fork34_outs_1_ready,
      clk => clk,
      rst => rst,
      outs => constant61_outs,
      outs_valid => constant61_outs_valid,
      outs_ready => constant61_outs_ready
    );

  extsi17 : entity work.extsi(arch) generic map(2, 32)
    port map(
      ins => constant61_outs,
      ins_valid => constant61_outs_valid,
      ins_ready => constant61_outs_ready,
      clk => clk,
      rst => rst,
      outs => extsi17_outs,
      outs_valid => extsi17_outs_valid,
      outs_ready => extsi17_outs_ready
    );

  constant62 : entity work.handshake_constant_0(arch) generic map(1)
    port map(
      ctrl_valid => fork34_outs_0_valid,
      ctrl_ready => fork34_outs_0_ready,
      clk => clk,
      rst => rst,
      outs => constant62_outs,
      outs_valid => constant62_outs_valid,
      outs_ready => constant62_outs_ready
    );

  fork35 : entity work.handshake_fork(arch) generic map(2, 1)
    port map(
      ins => constant62_outs,
      ins_valid => constant62_outs_valid,
      ins_ready => constant62_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork35_outs_0,
      outs(1) => fork35_outs_1,
      outs_valid(0) => fork35_outs_0_valid,
      outs_valid(1) => fork35_outs_1_valid,
      outs_ready(0) => fork35_outs_0_ready,
      outs_ready(1) => fork35_outs_1_ready
    );

  extsi19 : entity work.extsi(arch) generic map(1, 32)
    port map(
      ins => fork35_outs_1,
      ins_valid => fork35_outs_1_valid,
      ins_ready => fork35_outs_1_ready,
      clk => clk,
      rst => rst,
      outs => extsi19_outs,
      outs_valid => extsi19_outs_valid,
      outs_ready => extsi19_outs_ready
    );

  source9 : entity work.source(arch)
    port map(
      clk => clk,
      rst => rst,
      outs_valid => source9_outs_valid,
      outs_ready => source9_outs_ready
    );

  constant63 : entity work.handshake_constant_1(arch) generic map(2)
    port map(
      ctrl_valid => source9_outs_valid,
      ctrl_ready => source9_outs_ready,
      clk => clk,
      rst => rst,
      outs => constant63_outs,
      outs_valid => constant63_outs_valid,
      outs_ready => constant63_outs_ready
    );

  extsi20 : entity work.extsi(arch) generic map(2, 32)
    port map(
      ins => constant63_outs,
      ins_valid => constant63_outs_valid,
      ins_ready => constant63_outs_ready,
      clk => clk,
      rst => rst,
      outs => extsi20_outs,
      outs_valid => extsi20_outs_valid,
      outs_ready => extsi20_outs_ready
    );

  source10 : entity work.source(arch)
    port map(
      clk => clk,
      rst => rst,
      outs_valid => source10_outs_valid,
      outs_ready => source10_outs_ready
    );

  constant64 : entity work.handshake_constant_2(arch) generic map(3)
    port map(
      ctrl_valid => source10_outs_valid,
      ctrl_ready => source10_outs_ready,
      clk => clk,
      rst => rst,
      outs => constant64_outs,
      outs_valid => constant64_outs_valid,
      outs_ready => constant64_outs_ready
    );

  extsi21 : entity work.extsi(arch) generic map(3, 32)
    port map(
      ins => constant64_outs,
      ins_valid => constant64_outs_valid,
      ins_ready => constant64_outs_ready,
      clk => clk,
      rst => rst,
      outs => extsi21_outs,
      outs_valid => extsi21_outs_valid,
      outs_ready => extsi21_outs_ready
    );

  shli10 : entity work.shli(arch) generic map(32)
    port map(
      lhs => fork32_outs_0,
      lhs_valid => fork32_outs_0_valid,
      lhs_ready => fork32_outs_0_ready,
      rhs => extsi20_outs,
      rhs_valid => extsi20_outs_valid,
      rhs_ready => extsi20_outs_ready,
      clk => clk,
      rst => rst,
      result => shli10_result,
      result_valid => shli10_result_valid,
      result_ready => shli10_result_ready
    );

  buffer81 : entity work.oehb(arch) generic map(32)
    port map(
      ins => shli10_result,
      ins_valid => shli10_result_valid,
      ins_ready => shli10_result_ready,
      clk => clk,
      rst => rst,
      outs => buffer81_outs,
      outs_valid => buffer81_outs_valid,
      outs_ready => buffer81_outs_ready
    );

  trunci11 : entity work.trunci(arch) generic map(32, 7)
    port map(
      ins => buffer81_outs,
      ins_valid => buffer81_outs_valid,
      ins_ready => buffer81_outs_ready,
      clk => clk,
      rst => rst,
      outs => trunci11_outs,
      outs_valid => trunci11_outs_valid,
      outs_ready => trunci11_outs_ready
    );

  shli11 : entity work.shli(arch) generic map(32)
    port map(
      lhs => fork32_outs_1,
      lhs_valid => fork32_outs_1_valid,
      lhs_ready => fork32_outs_1_ready,
      rhs => extsi21_outs,
      rhs_valid => extsi21_outs_valid,
      rhs_ready => extsi21_outs_ready,
      clk => clk,
      rst => rst,
      result => shli11_result,
      result_valid => shli11_result_valid,
      result_ready => shli11_result_ready
    );

  buffer82 : entity work.oehb(arch) generic map(32)
    port map(
      ins => shli11_result,
      ins_valid => shli11_result_valid,
      ins_ready => shli11_result_ready,
      clk => clk,
      rst => rst,
      outs => buffer82_outs,
      outs_valid => buffer82_outs_valid,
      outs_ready => buffer82_outs_ready
    );

  trunci12 : entity work.trunci(arch) generic map(32, 7)
    port map(
      ins => buffer82_outs,
      ins_valid => buffer82_outs_valid,
      ins_ready => buffer82_outs_ready,
      clk => clk,
      rst => rst,
      outs => trunci12_outs,
      outs_valid => trunci12_outs_valid,
      outs_ready => trunci12_outs_ready
    );

  addi32 : entity work.addi(arch) generic map(7)
    port map(
      lhs => trunci11_outs,
      lhs_valid => trunci11_outs_valid,
      lhs_ready => trunci11_outs_ready,
      rhs => trunci12_outs,
      rhs_valid => trunci12_outs_valid,
      rhs_ready => trunci12_outs_ready,
      clk => clk,
      rst => rst,
      result => addi32_result,
      result_valid => addi32_result_valid,
      result_ready => addi32_result_ready
    );

  buffer83 : entity work.oehb(arch) generic map(7)
    port map(
      ins => addi32_result,
      ins_valid => addi32_result_valid,
      ins_ready => addi32_result_ready,
      clk => clk,
      rst => rst,
      outs => buffer83_outs,
      outs_valid => buffer83_outs_valid,
      outs_ready => buffer83_outs_ready
    );

  addi8 : entity work.addi(arch) generic map(7)
    port map(
      lhs => extsi70_outs,
      lhs_valid => extsi70_outs_valid,
      lhs_ready => extsi70_outs_ready,
      rhs => buffer83_outs,
      rhs_valid => buffer83_outs_valid,
      rhs_ready => buffer83_outs_ready,
      clk => clk,
      rst => rst,
      result => addi8_result,
      result_valid => addi8_result_valid,
      result_ready => addi8_result_ready
    );

  buffer2 : entity work.tfifo_dataless(arch) generic map(1)
    port map(
      ins_valid => store2_doneOut_valid,
      ins_ready => store2_doneOut_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer2_outs_valid,
      outs_ready => buffer2_outs_ready
    );

  fork36 : entity work.fork_dataless(arch) generic map(2)
    port map(
      ins_valid => buffer2_outs_valid,
      ins_ready => buffer2_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid(0) => fork36_outs_0_valid,
      outs_valid(1) => fork36_outs_1_valid,
      outs_ready(0) => fork36_outs_0_ready,
      outs_ready(1) => fork36_outs_1_ready
    );

  buffer84 : entity work.oehb(arch) generic map(7)
    port map(
      ins => addi8_result,
      ins_valid => addi8_result_valid,
      ins_ready => addi8_result_ready,
      clk => clk,
      rst => rst,
      outs => buffer84_outs,
      outs_valid => buffer84_outs_valid,
      outs_ready => buffer84_outs_ready
    );

  store2 : entity work.store(arch) generic map(32, 7)
    port map(
      addrIn => buffer84_outs,
      addrIn_valid => buffer84_outs_valid,
      addrIn_ready => buffer84_outs_ready,
      dataIn => extsi19_outs,
      dataIn_valid => extsi19_outs_valid,
      dataIn_ready => extsi19_outs_ready,
      doneFromMem_valid => mem_controller5_stDone_0_valid,
      doneFromMem_ready => mem_controller5_stDone_0_ready,
      clk => clk,
      rst => rst,
      addrOut => store2_addrOut,
      addrOut_valid => store2_addrOut_valid,
      addrOut_ready => store2_addrOut_ready,
      dataToMem => store2_dataToMem,
      dataToMem_valid => store2_dataToMem_valid,
      dataToMem_ready => store2_dataToMem_ready,
      doneOut_valid => store2_doneOut_valid,
      doneOut_ready => store2_doneOut_ready
    );

  extsi48 : entity work.extsi(arch) generic map(1, 5)
    port map(
      ins => fork35_outs_0,
      ins_valid => fork35_outs_0_valid,
      ins_ready => fork35_outs_0_ready,
      clk => clk,
      rst => rst,
      outs => extsi48_outs,
      outs_valid => extsi48_outs_valid,
      outs_ready => extsi48_outs_ready
    );

  cond_br122 : entity work.cond_br_dataless(arch)
    port map(
      condition => buffer86_outs,
      condition_valid => buffer86_outs_valid,
      condition_ready => buffer86_outs_ready,
      data_valid => fork38_outs_2_valid,
      data_ready => fork38_outs_2_ready,
      clk => clk,
      rst => rst,
      trueOut_valid => cond_br122_trueOut_valid,
      trueOut_ready => cond_br122_trueOut_ready,
      falseOut_valid => cond_br122_falseOut_valid,
      falseOut_ready => cond_br122_falseOut_ready
    );

  buffer86 : entity work.tfifo(arch) generic map(2, 1)
    port map(
      ins => fork51_outs_5,
      ins_valid => fork51_outs_5_valid,
      ins_ready => fork51_outs_5_ready,
      clk => clk,
      rst => rst,
      outs => buffer86_outs,
      outs_valid => buffer86_outs_valid,
      outs_ready => buffer86_outs_ready
    );

  sink9 : entity work.sink_dataless(arch)
    port map(
      ins_valid => cond_br122_falseOut_valid,
      ins_ready => cond_br122_falseOut_ready,
      clk => clk,
      rst => rst
    );

  buffer126 : entity work.oehb_dataless(arch)
    port map(
      ins_valid => buffer3_outs_valid,
      ins_ready => buffer3_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer126_outs_valid,
      outs_ready => buffer126_outs_ready
    );

  cond_br123 : entity work.cond_br_dataless(arch)
    port map(
      condition => buffer87_outs,
      condition_valid => buffer87_outs_valid,
      condition_ready => buffer87_outs_ready,
      data_valid => buffer126_outs_valid,
      data_ready => buffer126_outs_ready,
      clk => clk,
      rst => rst,
      trueOut_valid => cond_br123_trueOut_valid,
      trueOut_ready => cond_br123_trueOut_ready,
      falseOut_valid => cond_br123_falseOut_valid,
      falseOut_ready => cond_br123_falseOut_ready
    );

  buffer87 : entity work.tfifo(arch) generic map(3, 1)
    port map(
      ins => fork51_outs_4,
      ins_valid => fork51_outs_4_valid,
      ins_ready => fork51_outs_4_ready,
      clk => clk,
      rst => rst,
      outs => buffer87_outs,
      outs_valid => buffer87_outs_valid,
      outs_ready => buffer87_outs_ready
    );

  init24 : entity work.tehb_init(arch) generic map(1, 0)
    port map(
      ins => fork51_outs_3,
      ins_valid => fork51_outs_3_valid,
      ins_ready => fork51_outs_3_ready,
      clk => clk,
      rst => rst,
      outs => init24_outs,
      outs_valid => init24_outs_valid,
      outs_ready => init24_outs_ready
    );

  fork37 : entity work.handshake_fork(arch) generic map(2, 1)
    port map(
      ins => init24_outs,
      ins_valid => init24_outs_valid,
      ins_ready => init24_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork37_outs_0,
      outs(1) => fork37_outs_1,
      outs_valid(0) => fork37_outs_0_valid,
      outs_valid(1) => fork37_outs_1_valid,
      outs_ready(0) => fork37_outs_0_ready,
      outs_ready(1) => fork37_outs_1_ready
    );

  mux42 : entity work.mux_dataless(arch) generic map(2, 1)
    port map(
      index => buffer89_outs,
      index_valid => buffer89_outs_valid,
      index_ready => buffer89_outs_ready,
      ins_valid(0) => fork36_outs_1_valid,
      ins_valid(1) => cond_br122_trueOut_valid,
      ins_ready(0) => fork36_outs_1_ready,
      ins_ready(1) => cond_br122_trueOut_ready,
      clk => clk,
      rst => rst,
      outs_valid => mux42_outs_valid,
      outs_ready => mux42_outs_ready
    );

  buffer89 : entity work.tfifo(arch) generic map(2, 1)
    port map(
      ins => fork37_outs_1,
      ins_valid => fork37_outs_1_valid,
      ins_ready => fork37_outs_1_ready,
      clk => clk,
      rst => rst,
      outs => buffer89_outs,
      outs_valid => buffer89_outs_valid,
      outs_ready => buffer89_outs_ready
    );

  buffer85 : entity work.oehb_dataless(arch)
    port map(
      ins_valid => mux42_outs_valid,
      ins_ready => mux42_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer85_outs_valid,
      outs_ready => buffer85_outs_ready
    );

  buffer88 : entity work.tehb_dataless(arch)
    port map(
      ins_valid => buffer85_outs_valid,
      ins_ready => buffer85_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer88_outs_valid,
      outs_ready => buffer88_outs_ready
    );

  fork38 : entity work.fork_dataless(arch) generic map(3)
    port map(
      ins_valid => buffer88_outs_valid,
      ins_ready => buffer88_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid(0) => fork38_outs_0_valid,
      outs_valid(1) => fork38_outs_1_valid,
      outs_valid(2) => fork38_outs_2_valid,
      outs_ready(0) => fork38_outs_0_ready,
      outs_ready(1) => fork38_outs_1_ready,
      outs_ready(2) => fork38_outs_2_ready
    );

  buffer76 : entity work.oehb_dataless(arch)
    port map(
      ins_valid => mux40_outs_valid,
      ins_ready => mux40_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer76_outs_valid,
      outs_ready => buffer76_outs_ready
    );

  buffer77 : entity work.tehb_dataless(arch)
    port map(
      ins_valid => buffer76_outs_valid,
      ins_ready => buffer76_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer77_outs_valid,
      outs_ready => buffer77_outs_ready
    );

  mux45 : entity work.mux_dataless(arch) generic map(2, 1)
    port map(
      index => buffer90_outs,
      index_valid => buffer90_outs_valid,
      index_ready => buffer90_outs_ready,
      ins_valid(0) => buffer77_outs_valid,
      ins_valid(1) => cond_br123_trueOut_valid,
      ins_ready(0) => buffer77_outs_ready,
      ins_ready(1) => cond_br123_trueOut_ready,
      clk => clk,
      rst => rst,
      outs_valid => mux45_outs_valid,
      outs_ready => mux45_outs_ready
    );

  buffer90 : entity work.tfifo(arch) generic map(3, 1)
    port map(
      ins => fork37_outs_0,
      ins_valid => fork37_outs_0_valid,
      ins_ready => fork37_outs_0_ready,
      clk => clk,
      rst => rst,
      outs => buffer90_outs,
      outs_valid => buffer90_outs_valid,
      outs_ready => buffer90_outs_ready
    );

  mux9 : entity work.mux(arch) generic map(2, 5, 1)
    port map(
      index => fork45_outs_2,
      index_valid => fork45_outs_2_valid,
      index_ready => fork45_outs_2_ready,
      ins(0) => extsi48_outs,
      ins(1) => cond_br19_trueOut,
      ins_valid(0) => extsi48_outs_valid,
      ins_valid(1) => cond_br19_trueOut_valid,
      ins_ready(0) => extsi48_outs_ready,
      ins_ready(1) => cond_br19_trueOut_ready,
      clk => clk,
      rst => rst,
      outs => mux9_outs,
      outs_valid => mux9_outs_valid,
      outs_ready => mux9_outs_ready
    );

  buffer92 : entity work.oehb(arch) generic map(5)
    port map(
      ins => mux9_outs,
      ins_valid => mux9_outs_valid,
      ins_ready => mux9_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer92_outs,
      outs_valid => buffer92_outs_valid,
      outs_ready => buffer92_outs_ready
    );

  buffer93 : entity work.tehb(arch) generic map(5)
    port map(
      ins => buffer92_outs,
      ins_valid => buffer92_outs_valid,
      ins_ready => buffer92_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer93_outs,
      outs_valid => buffer93_outs_valid,
      outs_ready => buffer93_outs_ready
    );

  fork39 : entity work.handshake_fork(arch) generic map(3, 5)
    port map(
      ins => buffer93_outs,
      ins_valid => buffer93_outs_valid,
      ins_ready => buffer93_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork39_outs_0,
      outs(1) => fork39_outs_1,
      outs(2) => fork39_outs_2,
      outs_valid(0) => fork39_outs_0_valid,
      outs_valid(1) => fork39_outs_1_valid,
      outs_valid(2) => fork39_outs_2_valid,
      outs_ready(0) => fork39_outs_0_ready,
      outs_ready(1) => fork39_outs_1_ready,
      outs_ready(2) => fork39_outs_2_ready
    );

  extsi72 : entity work.extsi(arch) generic map(5, 7)
    port map(
      ins => fork39_outs_0,
      ins_valid => fork39_outs_0_valid,
      ins_ready => fork39_outs_0_ready,
      clk => clk,
      rst => rst,
      outs => extsi72_outs,
      outs_valid => extsi72_outs_valid,
      outs_ready => extsi72_outs_ready
    );

  extsi73 : entity work.extsi(arch) generic map(5, 6)
    port map(
      ins => fork39_outs_1,
      ins_valid => fork39_outs_1_valid,
      ins_ready => fork39_outs_1_ready,
      clk => clk,
      rst => rst,
      outs => extsi73_outs,
      outs_valid => extsi73_outs_valid,
      outs_ready => extsi73_outs_ready
    );

  extsi74 : entity work.extsi(arch) generic map(5, 32)
    port map(
      ins => fork39_outs_2,
      ins_valid => fork39_outs_2_valid,
      ins_ready => fork39_outs_2_ready,
      clk => clk,
      rst => rst,
      outs => extsi74_outs,
      outs_valid => extsi74_outs_valid,
      outs_ready => extsi74_outs_ready
    );

  fork40 : entity work.handshake_fork(arch) generic map(2, 32)
    port map(
      ins => extsi74_outs,
      ins_valid => extsi74_outs_valid,
      ins_ready => extsi74_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork40_outs_0,
      outs(1) => fork40_outs_1,
      outs_valid(0) => fork40_outs_0_valid,
      outs_valid(1) => fork40_outs_1_valid,
      outs_ready(0) => fork40_outs_0_ready,
      outs_ready(1) => fork40_outs_1_ready
    );

  mux10 : entity work.mux(arch) generic map(2, 5, 1)
    port map(
      index => fork45_outs_0,
      index_valid => fork45_outs_0_valid,
      index_ready => fork45_outs_0_ready,
      ins(0) => fork31_outs_0,
      ins(1) => cond_br20_trueOut,
      ins_valid(0) => fork31_outs_0_valid,
      ins_valid(1) => cond_br20_trueOut_valid,
      ins_ready(0) => fork31_outs_0_ready,
      ins_ready(1) => cond_br20_trueOut_ready,
      clk => clk,
      rst => rst,
      outs => mux10_outs,
      outs_valid => mux10_outs_valid,
      outs_ready => mux10_outs_ready
    );

  buffer94 : entity work.oehb(arch) generic map(5)
    port map(
      ins => mux10_outs,
      ins_valid => mux10_outs_valid,
      ins_ready => mux10_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer94_outs,
      outs_valid => buffer94_outs_valid,
      outs_ready => buffer94_outs_ready
    );

  buffer95 : entity work.tehb(arch) generic map(5)
    port map(
      ins => buffer94_outs,
      ins_valid => buffer94_outs_valid,
      ins_ready => buffer94_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer95_outs,
      outs_valid => buffer95_outs_valid,
      outs_ready => buffer95_outs_ready
    );

  fork41 : entity work.handshake_fork(arch) generic map(2, 5)
    port map(
      ins => buffer95_outs,
      ins_valid => buffer95_outs_valid,
      ins_ready => buffer95_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork41_outs_0,
      outs(1) => fork41_outs_1,
      outs_valid(0) => fork41_outs_0_valid,
      outs_valid(1) => fork41_outs_1_valid,
      outs_ready(0) => fork41_outs_0_ready,
      outs_ready(1) => fork41_outs_1_ready
    );

  extsi75 : entity work.extsi(arch) generic map(5, 32)
    port map(
      ins => fork41_outs_1,
      ins_valid => fork41_outs_1_valid,
      ins_ready => fork41_outs_1_ready,
      clk => clk,
      rst => rst,
      outs => extsi75_outs,
      outs_valid => extsi75_outs_valid,
      outs_ready => extsi75_outs_ready
    );

  fork42 : entity work.handshake_fork(arch) generic map(6, 32)
    port map(
      ins => extsi75_outs,
      ins_valid => extsi75_outs_valid,
      ins_ready => extsi75_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork42_outs_0,
      outs(1) => fork42_outs_1,
      outs(2) => fork42_outs_2,
      outs(3) => fork42_outs_3,
      outs(4) => fork42_outs_4,
      outs(5) => fork42_outs_5,
      outs_valid(0) => fork42_outs_0_valid,
      outs_valid(1) => fork42_outs_1_valid,
      outs_valid(2) => fork42_outs_2_valid,
      outs_valid(3) => fork42_outs_3_valid,
      outs_valid(4) => fork42_outs_4_valid,
      outs_valid(5) => fork42_outs_5_valid,
      outs_ready(0) => fork42_outs_0_ready,
      outs_ready(1) => fork42_outs_1_ready,
      outs_ready(2) => fork42_outs_2_ready,
      outs_ready(3) => fork42_outs_3_ready,
      outs_ready(4) => fork42_outs_4_ready,
      outs_ready(5) => fork42_outs_5_ready
    );

  mux11 : entity work.mux(arch) generic map(2, 5, 1)
    port map(
      index => buffer97_outs,
      index_valid => buffer97_outs_valid,
      index_ready => buffer97_outs_ready,
      ins(0) => fork30_outs_1,
      ins(1) => cond_br21_trueOut,
      ins_valid(0) => fork30_outs_1_valid,
      ins_valid(1) => cond_br21_trueOut_valid,
      ins_ready(0) => fork30_outs_1_ready,
      ins_ready(1) => cond_br21_trueOut_ready,
      clk => clk,
      rst => rst,
      outs => mux11_outs,
      outs_valid => mux11_outs_valid,
      outs_ready => mux11_outs_ready
    );

  buffer97 : entity work.tfifo(arch) generic map(1, 1)
    port map(
      ins => fork45_outs_1,
      ins_valid => fork45_outs_1_valid,
      ins_ready => fork45_outs_1_ready,
      clk => clk,
      rst => rst,
      outs => buffer97_outs,
      outs_valid => buffer97_outs_valid,
      outs_ready => buffer97_outs_ready
    );

  buffer96 : entity work.oehb(arch) generic map(5)
    port map(
      ins => mux11_outs,
      ins_valid => mux11_outs_valid,
      ins_ready => mux11_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer96_outs,
      outs_valid => buffer96_outs_valid,
      outs_ready => buffer96_outs_ready
    );

  buffer98 : entity work.tehb(arch) generic map(5)
    port map(
      ins => buffer96_outs,
      ins_valid => buffer96_outs_valid,
      ins_ready => buffer96_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer98_outs,
      outs_valid => buffer98_outs_valid,
      outs_ready => buffer98_outs_ready
    );

  fork43 : entity work.handshake_fork(arch) generic map(3, 5)
    port map(
      ins => buffer98_outs,
      ins_valid => buffer98_outs_valid,
      ins_ready => buffer98_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork43_outs_0,
      outs(1) => fork43_outs_1,
      outs(2) => fork43_outs_2,
      outs_valid(0) => fork43_outs_0_valid,
      outs_valid(1) => fork43_outs_1_valid,
      outs_valid(2) => fork43_outs_2_valid,
      outs_ready(0) => fork43_outs_0_ready,
      outs_ready(1) => fork43_outs_1_ready,
      outs_ready(2) => fork43_outs_2_ready
    );

  extsi76 : entity work.extsi(arch) generic map(5, 7)
    port map(
      ins => fork43_outs_0,
      ins_valid => fork43_outs_0_valid,
      ins_ready => fork43_outs_0_ready,
      clk => clk,
      rst => rst,
      outs => extsi76_outs,
      outs_valid => extsi76_outs_valid,
      outs_ready => extsi76_outs_ready
    );

  extsi77 : entity work.extsi(arch) generic map(5, 32)
    port map(
      ins => buffer99_outs,
      ins_valid => buffer99_outs_valid,
      ins_ready => buffer99_outs_ready,
      clk => clk,
      rst => rst,
      outs => extsi77_outs,
      outs_valid => extsi77_outs_valid,
      outs_ready => extsi77_outs_ready
    );

  buffer99 : entity work.tfifo(arch) generic map(3, 5)
    port map(
      ins => fork43_outs_2,
      ins_valid => fork43_outs_2_valid,
      ins_ready => fork43_outs_2_ready,
      clk => clk,
      rst => rst,
      outs => buffer99_outs,
      outs_valid => buffer99_outs_valid,
      outs_ready => buffer99_outs_ready
    );

  fork44 : entity work.handshake_fork(arch) generic map(2, 32)
    port map(
      ins => extsi77_outs,
      ins_valid => extsi77_outs_valid,
      ins_ready => extsi77_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork44_outs_0,
      outs(1) => fork44_outs_1,
      outs_valid(0) => fork44_outs_0_valid,
      outs_valid(1) => fork44_outs_1_valid,
      outs_ready(0) => fork44_outs_0_ready,
      outs_ready(1) => fork44_outs_1_ready
    );

  control_merge7 : entity work.control_merge_dataless(arch) generic map(2, 1)
    port map(
      ins_valid(0) => fork34_outs_2_valid,
      ins_valid(1) => cond_br22_trueOut_valid,
      ins_ready(0) => fork34_outs_2_ready,
      ins_ready(1) => cond_br22_trueOut_ready,
      clk => clk,
      rst => rst,
      outs_valid => control_merge7_outs_valid,
      outs_ready => control_merge7_outs_ready,
      index => control_merge7_index,
      index_valid => control_merge7_index_valid,
      index_ready => control_merge7_index_ready
    );

  fork45 : entity work.handshake_fork(arch) generic map(3, 1)
    port map(
      ins => control_merge7_index,
      ins_valid => control_merge7_index_valid,
      ins_ready => control_merge7_index_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork45_outs_0,
      outs(1) => fork45_outs_1,
      outs(2) => fork45_outs_2,
      outs_valid(0) => fork45_outs_0_valid,
      outs_valid(1) => fork45_outs_1_valid,
      outs_valid(2) => fork45_outs_2_valid,
      outs_ready(0) => fork45_outs_0_ready,
      outs_ready(1) => fork45_outs_1_ready,
      outs_ready(2) => fork45_outs_2_ready
    );

  buffer100 : entity work.oehb_dataless(arch)
    port map(
      ins_valid => control_merge7_outs_valid,
      ins_ready => control_merge7_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer100_outs_valid,
      outs_ready => buffer100_outs_ready
    );

  fork46 : entity work.fork_dataless(arch) generic map(2)
    port map(
      ins_valid => buffer100_outs_valid,
      ins_ready => buffer100_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid(0) => fork46_outs_0_valid,
      outs_valid(1) => fork46_outs_1_valid,
      outs_ready(0) => fork46_outs_0_ready,
      outs_ready(1) => fork46_outs_1_ready
    );

  constant65 : entity work.handshake_constant_1(arch) generic map(2)
    port map(
      ctrl_valid => fork46_outs_0_valid,
      ctrl_ready => fork46_outs_0_ready,
      clk => clk,
      rst => rst,
      outs => constant65_outs,
      outs_valid => constant65_outs_valid,
      outs_ready => constant65_outs_ready
    );

  extsi22 : entity work.extsi(arch) generic map(2, 32)
    port map(
      ins => constant65_outs,
      ins_valid => constant65_outs_valid,
      ins_ready => constant65_outs_ready,
      clk => clk,
      rst => rst,
      outs => extsi22_outs,
      outs_valid => extsi22_outs_valid,
      outs_ready => extsi22_outs_ready
    );

  source11 : entity work.source(arch)
    port map(
      clk => clk,
      rst => rst,
      outs_valid => source11_outs_valid,
      outs_ready => source11_outs_ready
    );

  constant66 : entity work.handshake_constant_3(arch) generic map(5)
    port map(
      ctrl_valid => source11_outs_valid,
      ctrl_ready => source11_outs_ready,
      clk => clk,
      rst => rst,
      outs => constant66_outs,
      outs_valid => constant66_outs_valid,
      outs_ready => constant66_outs_ready
    );

  extsi78 : entity work.extsi(arch) generic map(5, 6)
    port map(
      ins => constant66_outs,
      ins_valid => constant66_outs_valid,
      ins_ready => constant66_outs_ready,
      clk => clk,
      rst => rst,
      outs => extsi78_outs,
      outs_valid => extsi78_outs_valid,
      outs_ready => extsi78_outs_ready
    );

  source12 : entity work.source(arch)
    port map(
      clk => clk,
      rst => rst,
      outs_valid => source12_outs_valid,
      outs_ready => source12_outs_ready
    );

  constant67 : entity work.handshake_constant_1(arch) generic map(2)
    port map(
      ctrl_valid => source12_outs_valid,
      ctrl_ready => source12_outs_ready,
      clk => clk,
      rst => rst,
      outs => constant67_outs,
      outs_valid => constant67_outs_valid,
      outs_ready => constant67_outs_ready
    );

  fork47 : entity work.handshake_fork(arch) generic map(2, 2)
    port map(
      ins => constant67_outs,
      ins_valid => constant67_outs_valid,
      ins_ready => constant67_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork47_outs_0,
      outs(1) => fork47_outs_1,
      outs_valid(0) => fork47_outs_0_valid,
      outs_valid(1) => fork47_outs_1_valid,
      outs_ready(0) => fork47_outs_0_ready,
      outs_ready(1) => fork47_outs_1_ready
    );

  extsi79 : entity work.extsi(arch) generic map(2, 6)
    port map(
      ins => fork47_outs_0,
      ins_valid => fork47_outs_0_valid,
      ins_ready => fork47_outs_0_ready,
      clk => clk,
      rst => rst,
      outs => extsi79_outs,
      outs_valid => extsi79_outs_valid,
      outs_ready => extsi79_outs_ready
    );

  extsi24 : entity work.extsi(arch) generic map(2, 32)
    port map(
      ins => fork47_outs_1,
      ins_valid => fork47_outs_1_valid,
      ins_ready => fork47_outs_1_ready,
      clk => clk,
      rst => rst,
      outs => extsi24_outs,
      outs_valid => extsi24_outs_valid,
      outs_ready => extsi24_outs_ready
    );

  fork48 : entity work.handshake_fork(arch) generic map(4, 32)
    port map(
      ins => extsi24_outs,
      ins_valid => extsi24_outs_valid,
      ins_ready => extsi24_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork48_outs_0,
      outs(1) => fork48_outs_1,
      outs(2) => fork48_outs_2,
      outs(3) => fork48_outs_3,
      outs_valid(0) => fork48_outs_0_valid,
      outs_valid(1) => fork48_outs_1_valid,
      outs_valid(2) => fork48_outs_2_valid,
      outs_valid(3) => fork48_outs_3_valid,
      outs_ready(0) => fork48_outs_0_ready,
      outs_ready(1) => fork48_outs_1_ready,
      outs_ready(2) => fork48_outs_2_ready,
      outs_ready(3) => fork48_outs_3_ready
    );

  source13 : entity work.source(arch)
    port map(
      clk => clk,
      rst => rst,
      outs_valid => source13_outs_valid,
      outs_ready => source13_outs_ready
    );

  constant68 : entity work.handshake_constant_2(arch) generic map(3)
    port map(
      ctrl_valid => source13_outs_valid,
      ctrl_ready => source13_outs_ready,
      clk => clk,
      rst => rst,
      outs => constant68_outs,
      outs_valid => constant68_outs_valid,
      outs_ready => constant68_outs_ready
    );

  extsi25 : entity work.extsi(arch) generic map(3, 32)
    port map(
      ins => constant68_outs,
      ins_valid => constant68_outs_valid,
      ins_ready => constant68_outs_ready,
      clk => clk,
      rst => rst,
      outs => extsi25_outs,
      outs_valid => extsi25_outs_valid,
      outs_ready => extsi25_outs_ready
    );

  fork49 : entity work.handshake_fork(arch) generic map(4, 32)
    port map(
      ins => extsi25_outs,
      ins_valid => extsi25_outs_valid,
      ins_ready => extsi25_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork49_outs_0,
      outs(1) => fork49_outs_1,
      outs(2) => fork49_outs_2,
      outs(3) => fork49_outs_3,
      outs_valid(0) => fork49_outs_0_valid,
      outs_valid(1) => fork49_outs_1_valid,
      outs_valid(2) => fork49_outs_2_valid,
      outs_valid(3) => fork49_outs_3_valid,
      outs_ready(0) => fork49_outs_0_ready,
      outs_ready(1) => fork49_outs_1_ready,
      outs_ready(2) => fork49_outs_2_ready,
      outs_ready(3) => fork49_outs_3_ready
    );

  shli12 : entity work.shli(arch) generic map(32)
    port map(
      lhs => buffer103_outs,
      lhs_valid => buffer103_outs_valid,
      lhs_ready => buffer103_outs_ready,
      rhs => fork48_outs_0,
      rhs_valid => fork48_outs_0_valid,
      rhs_ready => fork48_outs_0_ready,
      clk => clk,
      rst => rst,
      result => shli12_result,
      result_valid => shli12_result_valid,
      result_ready => shli12_result_ready
    );

  buffer103 : entity work.tfifo(arch) generic map(1, 32)
    port map(
      ins => fork42_outs_0,
      ins_valid => fork42_outs_0_valid,
      ins_ready => fork42_outs_0_ready,
      clk => clk,
      rst => rst,
      outs => buffer103_outs,
      outs_valid => buffer103_outs_valid,
      outs_ready => buffer103_outs_ready
    );

  buffer101 : entity work.oehb(arch) generic map(32)
    port map(
      ins => shli12_result,
      ins_valid => shli12_result_valid,
      ins_ready => shli12_result_ready,
      clk => clk,
      rst => rst,
      outs => buffer101_outs,
      outs_valid => buffer101_outs_valid,
      outs_ready => buffer101_outs_ready
    );

  trunci13 : entity work.trunci(arch) generic map(32, 7)
    port map(
      ins => buffer101_outs,
      ins_valid => buffer101_outs_valid,
      ins_ready => buffer101_outs_ready,
      clk => clk,
      rst => rst,
      outs => trunci13_outs,
      outs_valid => trunci13_outs_valid,
      outs_ready => trunci13_outs_ready
    );

  shli13 : entity work.shli(arch) generic map(32)
    port map(
      lhs => buffer105_outs,
      lhs_valid => buffer105_outs_valid,
      lhs_ready => buffer105_outs_ready,
      rhs => fork49_outs_0,
      rhs_valid => fork49_outs_0_valid,
      rhs_ready => fork49_outs_0_ready,
      clk => clk,
      rst => rst,
      result => shli13_result,
      result_valid => shli13_result_valid,
      result_ready => shli13_result_ready
    );

  buffer105 : entity work.tfifo(arch) generic map(1, 32)
    port map(
      ins => fork42_outs_1,
      ins_valid => fork42_outs_1_valid,
      ins_ready => fork42_outs_1_ready,
      clk => clk,
      rst => rst,
      outs => buffer105_outs,
      outs_valid => buffer105_outs_valid,
      outs_ready => buffer105_outs_ready
    );

  buffer102 : entity work.oehb(arch) generic map(32)
    port map(
      ins => shli13_result,
      ins_valid => shli13_result_valid,
      ins_ready => shli13_result_ready,
      clk => clk,
      rst => rst,
      outs => buffer102_outs,
      outs_valid => buffer102_outs_valid,
      outs_ready => buffer102_outs_ready
    );

  trunci14 : entity work.trunci(arch) generic map(32, 7)
    port map(
      ins => buffer102_outs,
      ins_valid => buffer102_outs_valid,
      ins_ready => buffer102_outs_ready,
      clk => clk,
      rst => rst,
      outs => trunci14_outs,
      outs_valid => trunci14_outs_valid,
      outs_ready => trunci14_outs_ready
    );

  addi33 : entity work.addi(arch) generic map(7)
    port map(
      lhs => trunci13_outs,
      lhs_valid => trunci13_outs_valid,
      lhs_ready => trunci13_outs_ready,
      rhs => trunci14_outs,
      rhs_valid => trunci14_outs_valid,
      rhs_ready => trunci14_outs_ready,
      clk => clk,
      rst => rst,
      result => addi33_result,
      result_valid => addi33_result_valid,
      result_ready => addi33_result_ready
    );

  buffer104 : entity work.oehb(arch) generic map(7)
    port map(
      ins => addi33_result,
      ins_valid => addi33_result_valid,
      ins_ready => addi33_result_ready,
      clk => clk,
      rst => rst,
      outs => buffer104_outs,
      outs_valid => buffer104_outs_valid,
      outs_ready => buffer104_outs_ready
    );

  addi9 : entity work.addi(arch) generic map(7)
    port map(
      lhs => extsi72_outs,
      lhs_valid => extsi72_outs_valid,
      lhs_ready => extsi72_outs_ready,
      rhs => buffer104_outs,
      rhs_valid => buffer104_outs_valid,
      rhs_ready => buffer104_outs_ready,
      clk => clk,
      rst => rst,
      result => addi9_result,
      result_valid => addi9_result_valid,
      result_ready => addi9_result_ready
    );

  load3 : entity work.load(arch) generic map(32, 7)
    port map(
      addrIn => addi9_result,
      addrIn_valid => addi9_result_valid,
      addrIn_ready => addi9_result_ready,
      dataFromMem => mem_controller8_ldData_0,
      dataFromMem_valid => mem_controller8_ldData_0_valid,
      dataFromMem_ready => mem_controller8_ldData_0_ready,
      clk => clk,
      rst => rst,
      addrOut => load3_addrOut,
      addrOut_valid => load3_addrOut_valid,
      addrOut_ready => load3_addrOut_ready,
      dataOut => load3_dataOut,
      dataOut_valid => load3_dataOut_valid,
      dataOut_ready => load3_dataOut_ready
    );

  shli14 : entity work.shli(arch) generic map(32)
    port map(
      lhs => buffer107_outs,
      lhs_valid => buffer107_outs_valid,
      lhs_ready => buffer107_outs_ready,
      rhs => fork48_outs_1,
      rhs_valid => fork48_outs_1_valid,
      rhs_ready => fork48_outs_1_ready,
      clk => clk,
      rst => rst,
      result => shli14_result,
      result_valid => shli14_result_valid,
      result_ready => shli14_result_ready
    );

  buffer107 : entity work.tfifo(arch) generic map(1, 32)
    port map(
      ins => fork40_outs_0,
      ins_valid => fork40_outs_0_valid,
      ins_ready => fork40_outs_0_ready,
      clk => clk,
      rst => rst,
      outs => buffer107_outs,
      outs_valid => buffer107_outs_valid,
      outs_ready => buffer107_outs_ready
    );

  buffer106 : entity work.oehb(arch) generic map(32)
    port map(
      ins => shli14_result,
      ins_valid => shli14_result_valid,
      ins_ready => shli14_result_ready,
      clk => clk,
      rst => rst,
      outs => buffer106_outs,
      outs_valid => buffer106_outs_valid,
      outs_ready => buffer106_outs_ready
    );

  trunci15 : entity work.trunci(arch) generic map(32, 7)
    port map(
      ins => buffer106_outs,
      ins_valid => buffer106_outs_valid,
      ins_ready => buffer106_outs_ready,
      clk => clk,
      rst => rst,
      outs => trunci15_outs,
      outs_valid => trunci15_outs_valid,
      outs_ready => trunci15_outs_ready
    );

  shli15 : entity work.shli(arch) generic map(32)
    port map(
      lhs => buffer109_outs,
      lhs_valid => buffer109_outs_valid,
      lhs_ready => buffer109_outs_ready,
      rhs => fork49_outs_1,
      rhs_valid => fork49_outs_1_valid,
      rhs_ready => fork49_outs_1_ready,
      clk => clk,
      rst => rst,
      result => shli15_result,
      result_valid => shli15_result_valid,
      result_ready => shli15_result_ready
    );

  buffer109 : entity work.tfifo(arch) generic map(1, 32)
    port map(
      ins => fork40_outs_1,
      ins_valid => fork40_outs_1_valid,
      ins_ready => fork40_outs_1_ready,
      clk => clk,
      rst => rst,
      outs => buffer109_outs,
      outs_valid => buffer109_outs_valid,
      outs_ready => buffer109_outs_ready
    );

  buffer108 : entity work.oehb(arch) generic map(32)
    port map(
      ins => shli15_result,
      ins_valid => shli15_result_valid,
      ins_ready => shli15_result_ready,
      clk => clk,
      rst => rst,
      outs => buffer108_outs,
      outs_valid => buffer108_outs_valid,
      outs_ready => buffer108_outs_ready
    );

  trunci16 : entity work.trunci(arch) generic map(32, 7)
    port map(
      ins => buffer108_outs,
      ins_valid => buffer108_outs_valid,
      ins_ready => buffer108_outs_ready,
      clk => clk,
      rst => rst,
      outs => trunci16_outs,
      outs_valid => trunci16_outs_valid,
      outs_ready => trunci16_outs_ready
    );

  addi34 : entity work.addi(arch) generic map(7)
    port map(
      lhs => trunci15_outs,
      lhs_valid => trunci15_outs_valid,
      lhs_ready => trunci15_outs_ready,
      rhs => trunci16_outs,
      rhs_valid => trunci16_outs_valid,
      rhs_ready => trunci16_outs_ready,
      clk => clk,
      rst => rst,
      result => addi34_result,
      result_valid => addi34_result_valid,
      result_ready => addi34_result_ready
    );

  buffer114 : entity work.oehb(arch) generic map(7)
    port map(
      ins => addi34_result,
      ins_valid => addi34_result_valid,
      ins_ready => addi34_result_ready,
      clk => clk,
      rst => rst,
      outs => buffer114_outs,
      outs_valid => buffer114_outs_valid,
      outs_ready => buffer114_outs_ready
    );

  addi10 : entity work.addi(arch) generic map(7)
    port map(
      lhs => extsi76_outs,
      lhs_valid => extsi76_outs_valid,
      lhs_ready => extsi76_outs_ready,
      rhs => buffer114_outs,
      rhs_valid => buffer114_outs_valid,
      rhs_ready => buffer114_outs_ready,
      clk => clk,
      rst => rst,
      result => addi10_result,
      result_valid => addi10_result_valid,
      result_ready => addi10_result_ready
    );

  load4 : entity work.load(arch) generic map(32, 7)
    port map(
      addrIn => addi10_result,
      addrIn_valid => addi10_result_valid,
      addrIn_ready => addi10_result_ready,
      dataFromMem => mem_controller7_ldData_0,
      dataFromMem_valid => mem_controller7_ldData_0_valid,
      dataFromMem_ready => mem_controller7_ldData_0_ready,
      clk => clk,
      rst => rst,
      addrOut => load4_addrOut,
      addrOut_valid => load4_addrOut_valid,
      addrOut_ready => load4_addrOut_ready,
      dataOut => load4_dataOut,
      dataOut_valid => load4_dataOut_valid,
      dataOut_ready => load4_dataOut_ready
    );

  muli1 : entity work.muli(arch) generic map(32)
    port map(
      lhs => load3_dataOut,
      lhs_valid => load3_dataOut_valid,
      lhs_ready => load3_dataOut_ready,
      rhs => load4_dataOut,
      rhs_valid => load4_dataOut_valid,
      rhs_ready => load4_dataOut_ready,
      clk => clk,
      rst => rst,
      result => muli1_result,
      result_valid => muli1_result_valid,
      result_ready => muli1_result_ready
    );

  shli16 : entity work.shli(arch) generic map(32)
    port map(
      lhs => buffer111_outs,
      lhs_valid => buffer111_outs_valid,
      lhs_ready => buffer111_outs_ready,
      rhs => buffer110_outs,
      rhs_valid => buffer110_outs_valid,
      rhs_ready => buffer110_outs_ready,
      clk => clk,
      rst => rst,
      result => shli16_result,
      result_valid => shli16_result_valid,
      result_ready => shli16_result_ready
    );

  buffer110 : entity work.tfifo(arch) generic map(3, 32)
    port map(
      ins => fork48_outs_2,
      ins_valid => fork48_outs_2_valid,
      ins_ready => fork48_outs_2_ready,
      clk => clk,
      rst => rst,
      outs => buffer110_outs,
      outs_valid => buffer110_outs_valid,
      outs_ready => buffer110_outs_ready
    );

  buffer111 : entity work.tfifo(arch) generic map(2, 32)
    port map(
      ins => fork42_outs_2,
      ins_valid => fork42_outs_2_valid,
      ins_ready => fork42_outs_2_ready,
      clk => clk,
      rst => rst,
      outs => buffer111_outs,
      outs_valid => buffer111_outs_valid,
      outs_ready => buffer111_outs_ready
    );

  shli17 : entity work.shli(arch) generic map(32)
    port map(
      lhs => buffer113_outs,
      lhs_valid => buffer113_outs_valid,
      lhs_ready => buffer113_outs_ready,
      rhs => buffer112_outs,
      rhs_valid => buffer112_outs_valid,
      rhs_ready => buffer112_outs_ready,
      clk => clk,
      rst => rst,
      result => shli17_result,
      result_valid => shli17_result_valid,
      result_ready => shli17_result_ready
    );

  buffer112 : entity work.tfifo(arch) generic map(2, 32)
    port map(
      ins => fork49_outs_2,
      ins_valid => fork49_outs_2_valid,
      ins_ready => fork49_outs_2_ready,
      clk => clk,
      rst => rst,
      outs => buffer112_outs,
      outs_valid => buffer112_outs_valid,
      outs_ready => buffer112_outs_ready
    );

  buffer113 : entity work.tfifo(arch) generic map(2, 32)
    port map(
      ins => fork42_outs_3,
      ins_valid => fork42_outs_3_valid,
      ins_ready => fork42_outs_3_ready,
      clk => clk,
      rst => rst,
      outs => buffer113_outs,
      outs_valid => buffer113_outs_valid,
      outs_ready => buffer113_outs_ready
    );

  buffer119 : entity work.oehb(arch) generic map(32)
    port map(
      ins => shli16_result,
      ins_valid => shli16_result_valid,
      ins_ready => shli16_result_ready,
      clk => clk,
      rst => rst,
      outs => buffer119_outs,
      outs_valid => buffer119_outs_valid,
      outs_ready => buffer119_outs_ready
    );

  buffer120 : entity work.oehb(arch) generic map(32)
    port map(
      ins => shli17_result,
      ins_valid => shli17_result_valid,
      ins_ready => shli17_result_ready,
      clk => clk,
      rst => rst,
      outs => buffer120_outs,
      outs_valid => buffer120_outs_valid,
      outs_ready => buffer120_outs_ready
    );

  addi35 : entity work.addi(arch) generic map(32)
    port map(
      lhs => buffer119_outs,
      lhs_valid => buffer119_outs_valid,
      lhs_ready => buffer119_outs_ready,
      rhs => buffer120_outs,
      rhs_valid => buffer120_outs_valid,
      rhs_ready => buffer120_outs_ready,
      clk => clk,
      rst => rst,
      result => addi35_result,
      result_valid => addi35_result_valid,
      result_ready => addi35_result_ready
    );

  buffer122 : entity work.oehb(arch) generic map(32)
    port map(
      ins => addi35_result,
      ins_valid => addi35_result_valid,
      ins_ready => addi35_result_ready,
      clk => clk,
      rst => rst,
      outs => buffer122_outs,
      outs_valid => buffer122_outs_valid,
      outs_ready => buffer122_outs_ready
    );

  addi11 : entity work.addi(arch) generic map(32)
    port map(
      lhs => fork44_outs_0,
      lhs_valid => fork44_outs_0_valid,
      lhs_ready => fork44_outs_0_ready,
      rhs => buffer122_outs,
      rhs_valid => buffer122_outs_valid,
      rhs_ready => buffer122_outs_ready,
      clk => clk,
      rst => rst,
      result => addi11_result,
      result_valid => addi11_result_valid,
      result_ready => addi11_result_ready
    );

  buffer91 : entity work.tehb_dataless(arch)
    port map(
      ins_valid => mux45_outs_valid,
      ins_ready => mux45_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer91_outs_valid,
      outs_ready => buffer91_outs_ready
    );

  gate2 : entity work.gate(arch) generic map(3, 32)
    port map(
      ins(0) => addi11_result,
      ins_valid(0) => addi11_result_valid,
      ins_valid(1) => buffer91_outs_valid,
      ins_valid(2) => fork38_outs_1_valid,
      ins_ready(0) => addi11_result_ready,
      ins_ready(1) => buffer91_outs_ready,
      ins_ready(2) => fork38_outs_1_ready,
      clk => clk,
      rst => rst,
      outs => gate2_outs,
      outs_valid => gate2_outs_valid,
      outs_ready => gate2_outs_ready
    );

  trunci17 : entity work.trunci(arch) generic map(32, 7)
    port map(
      ins => gate2_outs,
      ins_valid => gate2_outs_valid,
      ins_ready => gate2_outs_ready,
      clk => clk,
      rst => rst,
      outs => trunci17_outs,
      outs_valid => trunci17_outs_valid,
      outs_ready => trunci17_outs_ready
    );

  load5 : entity work.load(arch) generic map(32, 7)
    port map(
      addrIn => trunci17_outs,
      addrIn_valid => trunci17_outs_valid,
      addrIn_ready => trunci17_outs_ready,
      dataFromMem => mem_controller5_ldData_0,
      dataFromMem_valid => mem_controller5_ldData_0_valid,
      dataFromMem_ready => mem_controller5_ldData_0_ready,
      clk => clk,
      rst => rst,
      addrOut => load5_addrOut,
      addrOut_valid => load5_addrOut_valid,
      addrOut_ready => load5_addrOut_ready,
      dataOut => load5_dataOut,
      dataOut_valid => load5_dataOut_valid,
      dataOut_ready => load5_dataOut_ready
    );

  addi1 : entity work.addi(arch) generic map(32)
    port map(
      lhs => load5_dataOut,
      lhs_valid => load5_dataOut_valid,
      lhs_ready => load5_dataOut_ready,
      rhs => muli1_result,
      rhs_valid => muli1_result_valid,
      rhs_ready => muli1_result_ready,
      clk => clk,
      rst => rst,
      result => addi1_result,
      result_valid => addi1_result_valid,
      result_ready => addi1_result_ready
    );

  shli18 : entity work.shli(arch) generic map(32)
    port map(
      lhs => buffer116_outs,
      lhs_valid => buffer116_outs_valid,
      lhs_ready => buffer116_outs_ready,
      rhs => buffer115_outs,
      rhs_valid => buffer115_outs_valid,
      rhs_ready => buffer115_outs_ready,
      clk => clk,
      rst => rst,
      result => shli18_result,
      result_valid => shli18_result_valid,
      result_ready => shli18_result_ready
    );

  buffer115 : entity work.tfifo(arch) generic map(3, 32)
    port map(
      ins => fork48_outs_3,
      ins_valid => fork48_outs_3_valid,
      ins_ready => fork48_outs_3_ready,
      clk => clk,
      rst => rst,
      outs => buffer115_outs,
      outs_valid => buffer115_outs_valid,
      outs_ready => buffer115_outs_ready
    );

  buffer116 : entity work.tfifo(arch) generic map(3, 32)
    port map(
      ins => fork42_outs_4,
      ins_valid => fork42_outs_4_valid,
      ins_ready => fork42_outs_4_ready,
      clk => clk,
      rst => rst,
      outs => buffer116_outs,
      outs_valid => buffer116_outs_valid,
      outs_ready => buffer116_outs_ready
    );

  shli19 : entity work.shli(arch) generic map(32)
    port map(
      lhs => buffer118_outs,
      lhs_valid => buffer118_outs_valid,
      lhs_ready => buffer118_outs_ready,
      rhs => buffer117_outs,
      rhs_valid => buffer117_outs_valid,
      rhs_ready => buffer117_outs_ready,
      clk => clk,
      rst => rst,
      result => shli19_result,
      result_valid => shli19_result_valid,
      result_ready => shli19_result_ready
    );

  buffer117 : entity work.tfifo(arch) generic map(3, 32)
    port map(
      ins => fork49_outs_3,
      ins_valid => fork49_outs_3_valid,
      ins_ready => fork49_outs_3_ready,
      clk => clk,
      rst => rst,
      outs => buffer117_outs,
      outs_valid => buffer117_outs_valid,
      outs_ready => buffer117_outs_ready
    );

  buffer118 : entity work.tfifo(arch) generic map(3, 32)
    port map(
      ins => fork42_outs_5,
      ins_valid => fork42_outs_5_valid,
      ins_ready => fork42_outs_5_ready,
      clk => clk,
      rst => rst,
      outs => buffer118_outs,
      outs_valid => buffer118_outs_valid,
      outs_ready => buffer118_outs_ready
    );

  buffer123 : entity work.oehb(arch) generic map(32)
    port map(
      ins => shli18_result,
      ins_valid => shli18_result_valid,
      ins_ready => shli18_result_ready,
      clk => clk,
      rst => rst,
      outs => buffer123_outs,
      outs_valid => buffer123_outs_valid,
      outs_ready => buffer123_outs_ready
    );

  buffer124 : entity work.oehb(arch) generic map(32)
    port map(
      ins => shli19_result,
      ins_valid => shli19_result_valid,
      ins_ready => shli19_result_ready,
      clk => clk,
      rst => rst,
      outs => buffer124_outs,
      outs_valid => buffer124_outs_valid,
      outs_ready => buffer124_outs_ready
    );

  addi36 : entity work.addi(arch) generic map(32)
    port map(
      lhs => buffer123_outs,
      lhs_valid => buffer123_outs_valid,
      lhs_ready => buffer123_outs_ready,
      rhs => buffer124_outs,
      rhs_valid => buffer124_outs_valid,
      rhs_ready => buffer124_outs_ready,
      clk => clk,
      rst => rst,
      result => addi36_result,
      result_valid => addi36_result_valid,
      result_ready => addi36_result_ready
    );

  buffer125 : entity work.oehb(arch) generic map(32)
    port map(
      ins => addi36_result,
      ins_valid => addi36_result_valid,
      ins_ready => addi36_result_ready,
      clk => clk,
      rst => rst,
      outs => buffer125_outs,
      outs_valid => buffer125_outs_valid,
      outs_ready => buffer125_outs_ready
    );

  addi12 : entity work.addi(arch) generic map(32)
    port map(
      lhs => fork44_outs_1,
      lhs_valid => fork44_outs_1_valid,
      lhs_ready => fork44_outs_1_ready,
      rhs => buffer125_outs,
      rhs_valid => buffer125_outs_valid,
      rhs_ready => buffer125_outs_ready,
      clk => clk,
      rst => rst,
      result => addi12_result,
      result_valid => addi12_result_valid,
      result_ready => addi12_result_ready
    );

  buffer3 : entity work.tfifo_dataless(arch) generic map(1)
    port map(
      ins_valid => store3_doneOut_valid,
      ins_ready => store3_doneOut_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer3_outs_valid,
      outs_ready => buffer3_outs_ready
    );

  gate3 : entity work.gate(arch) generic map(2, 32)
    port map(
      ins(0) => addi12_result,
      ins_valid(0) => addi12_result_valid,
      ins_valid(1) => fork38_outs_0_valid,
      ins_ready(0) => addi12_result_ready,
      ins_ready(1) => fork38_outs_0_ready,
      clk => clk,
      rst => rst,
      outs => gate3_outs,
      outs_valid => gate3_outs_valid,
      outs_ready => gate3_outs_ready
    );

  trunci18 : entity work.trunci(arch) generic map(32, 7)
    port map(
      ins => gate3_outs,
      ins_valid => gate3_outs_valid,
      ins_ready => gate3_outs_ready,
      clk => clk,
      rst => rst,
      outs => trunci18_outs,
      outs_valid => trunci18_outs_valid,
      outs_ready => trunci18_outs_ready
    );

  store3 : entity work.store(arch) generic map(32, 7)
    port map(
      addrIn => trunci18_outs,
      addrIn_valid => trunci18_outs_valid,
      addrIn_ready => trunci18_outs_ready,
      dataIn => addi1_result,
      dataIn_valid => addi1_result_valid,
      dataIn_ready => addi1_result_ready,
      doneFromMem_valid => mem_controller5_stDone_1_valid,
      doneFromMem_ready => mem_controller5_stDone_1_ready,
      clk => clk,
      rst => rst,
      addrOut => store3_addrOut,
      addrOut_valid => store3_addrOut_valid,
      addrOut_ready => store3_addrOut_ready,
      dataToMem => store3_dataToMem,
      dataToMem_valid => store3_dataToMem_valid,
      dataToMem_ready => store3_dataToMem_ready,
      doneOut_valid => store3_doneOut_valid,
      doneOut_ready => store3_doneOut_ready
    );

  addi21 : entity work.addi(arch) generic map(6)
    port map(
      lhs => extsi73_outs,
      lhs_valid => extsi73_outs_valid,
      lhs_ready => extsi73_outs_ready,
      rhs => extsi79_outs,
      rhs_valid => extsi79_outs_valid,
      rhs_ready => extsi79_outs_ready,
      clk => clk,
      rst => rst,
      result => addi21_result,
      result_valid => addi21_result_valid,
      result_ready => addi21_result_ready
    );

  fork50 : entity work.handshake_fork(arch) generic map(2, 6)
    port map(
      ins => addi21_result,
      ins_valid => addi21_result_valid,
      ins_ready => addi21_result_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork50_outs_0,
      outs(1) => fork50_outs_1,
      outs_valid(0) => fork50_outs_0_valid,
      outs_valid(1) => fork50_outs_1_valid,
      outs_ready(0) => fork50_outs_0_ready,
      outs_ready(1) => fork50_outs_1_ready
    );

  trunci19 : entity work.trunci(arch) generic map(6, 5)
    port map(
      ins => fork50_outs_0,
      ins_valid => fork50_outs_0_valid,
      ins_ready => fork50_outs_0_ready,
      clk => clk,
      rst => rst,
      outs => trunci19_outs,
      outs_valid => trunci19_outs_valid,
      outs_ready => trunci19_outs_ready
    );

  buffer131 : entity work.oehb(arch) generic map(6)
    port map(
      ins => buffer121_outs,
      ins_valid => buffer121_outs_valid,
      ins_ready => buffer121_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer131_outs,
      outs_valid => buffer131_outs_valid,
      outs_ready => buffer131_outs_ready
    );

  cmpi3 : entity work.handshake_cmpi_0(arch) generic map(6)
    port map(
      lhs => buffer131_outs,
      lhs_valid => buffer131_outs_valid,
      lhs_ready => buffer131_outs_ready,
      rhs => extsi78_outs,
      rhs_valid => extsi78_outs_valid,
      rhs_ready => extsi78_outs_ready,
      clk => clk,
      rst => rst,
      result => cmpi3_result,
      result_valid => cmpi3_result_valid,
      result_ready => cmpi3_result_ready
    );

  buffer121 : entity work.tfifo(arch) generic map(1, 6)
    port map(
      ins => fork50_outs_1,
      ins_valid => fork50_outs_1_valid,
      ins_ready => fork50_outs_1_ready,
      clk => clk,
      rst => rst,
      outs => buffer121_outs,
      outs_valid => buffer121_outs_valid,
      outs_ready => buffer121_outs_ready
    );

  buffer130 : entity work.oehb(arch) generic map(1)
    port map(
      ins => cmpi3_result,
      ins_valid => cmpi3_result_valid,
      ins_ready => cmpi3_result_ready,
      clk => clk,
      rst => rst,
      outs => buffer130_outs,
      outs_valid => buffer130_outs_valid,
      outs_ready => buffer130_outs_ready
    );

  fork51 : entity work.handshake_fork(arch) generic map(7, 1)
    port map(
      ins => buffer130_outs,
      ins_valid => buffer130_outs_valid,
      ins_ready => buffer130_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork51_outs_0,
      outs(1) => fork51_outs_1,
      outs(2) => fork51_outs_2,
      outs(3) => fork51_outs_3,
      outs(4) => fork51_outs_4,
      outs(5) => fork51_outs_5,
      outs(6) => fork51_outs_6,
      outs_valid(0) => fork51_outs_0_valid,
      outs_valid(1) => fork51_outs_1_valid,
      outs_valid(2) => fork51_outs_2_valid,
      outs_valid(3) => fork51_outs_3_valid,
      outs_valid(4) => fork51_outs_4_valid,
      outs_valid(5) => fork51_outs_5_valid,
      outs_valid(6) => fork51_outs_6_valid,
      outs_ready(0) => fork51_outs_0_ready,
      outs_ready(1) => fork51_outs_1_ready,
      outs_ready(2) => fork51_outs_2_ready,
      outs_ready(3) => fork51_outs_3_ready,
      outs_ready(4) => fork51_outs_4_ready,
      outs_ready(5) => fork51_outs_5_ready,
      outs_ready(6) => fork51_outs_6_ready
    );

  cond_br19 : entity work.cond_br(arch) generic map(5)
    port map(
      condition => fork51_outs_0,
      condition_valid => fork51_outs_0_valid,
      condition_ready => fork51_outs_0_ready,
      data => trunci19_outs,
      data_valid => trunci19_outs_valid,
      data_ready => trunci19_outs_ready,
      clk => clk,
      rst => rst,
      trueOut => cond_br19_trueOut,
      trueOut_valid => cond_br19_trueOut_valid,
      trueOut_ready => cond_br19_trueOut_ready,
      falseOut => cond_br19_falseOut,
      falseOut_valid => cond_br19_falseOut_valid,
      falseOut_ready => cond_br19_falseOut_ready
    );

  sink10 : entity work.sink(arch) generic map(5)
    port map(
      ins => cond_br19_falseOut,
      ins_valid => cond_br19_falseOut_valid,
      ins_ready => cond_br19_falseOut_ready,
      clk => clk,
      rst => rst
    );

  cond_br20 : entity work.cond_br(arch) generic map(5)
    port map(
      condition => fork51_outs_1,
      condition_valid => fork51_outs_1_valid,
      condition_ready => fork51_outs_1_ready,
      data => fork41_outs_0,
      data_valid => fork41_outs_0_valid,
      data_ready => fork41_outs_0_ready,
      clk => clk,
      rst => rst,
      trueOut => cond_br20_trueOut,
      trueOut_valid => cond_br20_trueOut_valid,
      trueOut_ready => cond_br20_trueOut_ready,
      falseOut => cond_br20_falseOut,
      falseOut_valid => cond_br20_falseOut_valid,
      falseOut_ready => cond_br20_falseOut_ready
    );

  cond_br21 : entity work.cond_br(arch) generic map(5)
    port map(
      condition => fork51_outs_2,
      condition_valid => fork51_outs_2_valid,
      condition_ready => fork51_outs_2_ready,
      data => fork43_outs_1,
      data_valid => fork43_outs_1_valid,
      data_ready => fork43_outs_1_ready,
      clk => clk,
      rst => rst,
      trueOut => cond_br21_trueOut,
      trueOut_valid => cond_br21_trueOut_valid,
      trueOut_ready => cond_br21_trueOut_ready,
      falseOut => cond_br21_falseOut,
      falseOut_valid => cond_br21_falseOut_valid,
      falseOut_ready => cond_br21_falseOut_ready
    );

  cond_br22 : entity work.cond_br_dataless(arch)
    port map(
      condition => buffer127_outs,
      condition_valid => buffer127_outs_valid,
      condition_ready => buffer127_outs_ready,
      data_valid => fork46_outs_1_valid,
      data_ready => fork46_outs_1_ready,
      clk => clk,
      rst => rst,
      trueOut_valid => cond_br22_trueOut_valid,
      trueOut_ready => cond_br22_trueOut_ready,
      falseOut_valid => cond_br22_falseOut_valid,
      falseOut_ready => cond_br22_falseOut_ready
    );

  buffer127 : entity work.tfifo(arch) generic map(1, 1)
    port map(
      ins => fork51_outs_6,
      ins_valid => fork51_outs_6_valid,
      ins_ready => fork51_outs_6_ready,
      clk => clk,
      rst => rst,
      outs => buffer127_outs,
      outs_valid => buffer127_outs_valid,
      outs_ready => buffer127_outs_ready
    );

  cond_br124 : entity work.cond_br_dataless(arch)
    port map(
      condition => buffer128_outs,
      condition_valid => buffer128_outs_valid,
      condition_ready => buffer128_outs_ready,
      data_valid => fork36_outs_0_valid,
      data_ready => fork36_outs_0_ready,
      clk => clk,
      rst => rst,
      trueOut_valid => cond_br124_trueOut_valid,
      trueOut_ready => cond_br124_trueOut_ready,
      falseOut_valid => cond_br124_falseOut_valid,
      falseOut_ready => cond_br124_falseOut_ready
    );

  buffer128 : entity work.tfifo(arch) generic map(1, 1)
    port map(
      ins => fork53_outs_3,
      ins_valid => fork53_outs_3_valid,
      ins_ready => fork53_outs_3_ready,
      clk => clk,
      rst => rst,
      outs => buffer128_outs,
      outs_valid => buffer128_outs_valid,
      outs_ready => buffer128_outs_ready
    );

  sink11 : entity work.sink_dataless(arch)
    port map(
      ins_valid => cond_br124_trueOut_valid,
      ins_ready => cond_br124_trueOut_ready,
      clk => clk,
      rst => rst
    );

  cond_br125 : entity work.cond_br_dataless(arch)
    port map(
      condition => buffer129_outs,
      condition_valid => buffer129_outs_valid,
      condition_ready => buffer129_outs_ready,
      data_valid => cond_br123_falseOut_valid,
      data_ready => cond_br123_falseOut_ready,
      clk => clk,
      rst => rst,
      trueOut_valid => cond_br125_trueOut_valid,
      trueOut_ready => cond_br125_trueOut_ready,
      falseOut_valid => cond_br125_falseOut_valid,
      falseOut_ready => cond_br125_falseOut_ready
    );

  buffer129 : entity work.tfifo(arch) generic map(1, 1)
    port map(
      ins => fork53_outs_2,
      ins_valid => fork53_outs_2_valid,
      ins_ready => fork53_outs_2_ready,
      clk => clk,
      rst => rst,
      outs => buffer129_outs,
      outs_valid => buffer129_outs_valid,
      outs_ready => buffer129_outs_ready
    );

  extsi80 : entity work.extsi(arch) generic map(5, 6)
    port map(
      ins => cond_br21_falseOut,
      ins_valid => cond_br21_falseOut_valid,
      ins_ready => cond_br21_falseOut_ready,
      clk => clk,
      rst => rst,
      outs => extsi80_outs,
      outs_valid => extsi80_outs_valid,
      outs_ready => extsi80_outs_ready
    );

  source14 : entity work.source(arch)
    port map(
      clk => clk,
      rst => rst,
      outs_valid => source14_outs_valid,
      outs_ready => source14_outs_ready
    );

  constant69 : entity work.handshake_constant_3(arch) generic map(5)
    port map(
      ctrl_valid => source14_outs_valid,
      ctrl_ready => source14_outs_ready,
      clk => clk,
      rst => rst,
      outs => constant69_outs,
      outs_valid => constant69_outs_valid,
      outs_ready => constant69_outs_ready
    );

  extsi81 : entity work.extsi(arch) generic map(5, 6)
    port map(
      ins => constant69_outs,
      ins_valid => constant69_outs_valid,
      ins_ready => constant69_outs_ready,
      clk => clk,
      rst => rst,
      outs => extsi81_outs,
      outs_valid => extsi81_outs_valid,
      outs_ready => extsi81_outs_ready
    );

  source15 : entity work.source(arch)
    port map(
      clk => clk,
      rst => rst,
      outs_valid => source15_outs_valid,
      outs_ready => source15_outs_ready
    );

  constant70 : entity work.handshake_constant_1(arch) generic map(2)
    port map(
      ctrl_valid => source15_outs_valid,
      ctrl_ready => source15_outs_ready,
      clk => clk,
      rst => rst,
      outs => constant70_outs,
      outs_valid => constant70_outs_valid,
      outs_ready => constant70_outs_ready
    );

  extsi82 : entity work.extsi(arch) generic map(2, 6)
    port map(
      ins => constant70_outs,
      ins_valid => constant70_outs_valid,
      ins_ready => constant70_outs_ready,
      clk => clk,
      rst => rst,
      outs => extsi82_outs,
      outs_valid => extsi82_outs_valid,
      outs_ready => extsi82_outs_ready
    );

  addi22 : entity work.addi(arch) generic map(6)
    port map(
      lhs => extsi80_outs,
      lhs_valid => extsi80_outs_valid,
      lhs_ready => extsi80_outs_ready,
      rhs => extsi82_outs,
      rhs_valid => extsi82_outs_valid,
      rhs_ready => extsi82_outs_ready,
      clk => clk,
      rst => rst,
      result => addi22_result,
      result_valid => addi22_result_valid,
      result_ready => addi22_result_ready
    );

  buffer132 : entity work.oehb(arch) generic map(6)
    port map(
      ins => addi22_result,
      ins_valid => addi22_result_valid,
      ins_ready => addi22_result_ready,
      clk => clk,
      rst => rst,
      outs => buffer132_outs,
      outs_valid => buffer132_outs_valid,
      outs_ready => buffer132_outs_ready
    );

  fork52 : entity work.handshake_fork(arch) generic map(2, 6)
    port map(
      ins => buffer132_outs,
      ins_valid => buffer132_outs_valid,
      ins_ready => buffer132_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork52_outs_0,
      outs(1) => fork52_outs_1,
      outs_valid(0) => fork52_outs_0_valid,
      outs_valid(1) => fork52_outs_1_valid,
      outs_ready(0) => fork52_outs_0_ready,
      outs_ready(1) => fork52_outs_1_ready
    );

  trunci20 : entity work.trunci(arch) generic map(6, 5)
    port map(
      ins => fork52_outs_0,
      ins_valid => fork52_outs_0_valid,
      ins_ready => fork52_outs_0_ready,
      clk => clk,
      rst => rst,
      outs => trunci20_outs,
      outs_valid => trunci20_outs_valid,
      outs_ready => trunci20_outs_ready
    );

  cmpi4 : entity work.handshake_cmpi_0(arch) generic map(6)
    port map(
      lhs => fork52_outs_1,
      lhs_valid => fork52_outs_1_valid,
      lhs_ready => fork52_outs_1_ready,
      rhs => extsi81_outs,
      rhs_valid => extsi81_outs_valid,
      rhs_ready => extsi81_outs_ready,
      clk => clk,
      rst => rst,
      result => cmpi4_result,
      result_valid => cmpi4_result_valid,
      result_ready => cmpi4_result_ready
    );

  buffer133 : entity work.oehb(arch) generic map(1)
    port map(
      ins => cmpi4_result,
      ins_valid => cmpi4_result_valid,
      ins_ready => cmpi4_result_ready,
      clk => clk,
      rst => rst,
      outs => buffer133_outs,
      outs_valid => buffer133_outs_valid,
      outs_ready => buffer133_outs_ready
    );

  fork53 : entity work.handshake_fork(arch) generic map(6, 1)
    port map(
      ins => buffer133_outs,
      ins_valid => buffer133_outs_valid,
      ins_ready => buffer133_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork53_outs_0,
      outs(1) => fork53_outs_1,
      outs(2) => fork53_outs_2,
      outs(3) => fork53_outs_3,
      outs(4) => fork53_outs_4,
      outs(5) => fork53_outs_5,
      outs_valid(0) => fork53_outs_0_valid,
      outs_valid(1) => fork53_outs_1_valid,
      outs_valid(2) => fork53_outs_2_valid,
      outs_valid(3) => fork53_outs_3_valid,
      outs_valid(4) => fork53_outs_4_valid,
      outs_valid(5) => fork53_outs_5_valid,
      outs_ready(0) => fork53_outs_0_ready,
      outs_ready(1) => fork53_outs_1_ready,
      outs_ready(2) => fork53_outs_2_ready,
      outs_ready(3) => fork53_outs_3_ready,
      outs_ready(4) => fork53_outs_4_ready,
      outs_ready(5) => fork53_outs_5_ready
    );

  cond_br23 : entity work.cond_br(arch) generic map(5)
    port map(
      condition => fork53_outs_0,
      condition_valid => fork53_outs_0_valid,
      condition_ready => fork53_outs_0_ready,
      data => trunci20_outs,
      data_valid => trunci20_outs_valid,
      data_ready => trunci20_outs_ready,
      clk => clk,
      rst => rst,
      trueOut => cond_br23_trueOut,
      trueOut_valid => cond_br23_trueOut_valid,
      trueOut_ready => cond_br23_trueOut_ready,
      falseOut => cond_br23_falseOut,
      falseOut_valid => cond_br23_falseOut_valid,
      falseOut_ready => cond_br23_falseOut_ready
    );

  sink13 : entity work.sink(arch) generic map(5)
    port map(
      ins => cond_br23_falseOut,
      ins_valid => cond_br23_falseOut_valid,
      ins_ready => cond_br23_falseOut_ready,
      clk => clk,
      rst => rst
    );

  cond_br24 : entity work.cond_br(arch) generic map(5)
    port map(
      condition => fork53_outs_1,
      condition_valid => fork53_outs_1_valid,
      condition_ready => fork53_outs_1_ready,
      data => cond_br20_falseOut,
      data_valid => cond_br20_falseOut_valid,
      data_ready => cond_br20_falseOut_ready,
      clk => clk,
      rst => rst,
      trueOut => cond_br24_trueOut,
      trueOut_valid => cond_br24_trueOut_valid,
      trueOut_ready => cond_br24_trueOut_ready,
      falseOut => cond_br24_falseOut,
      falseOut_valid => cond_br24_falseOut_valid,
      falseOut_ready => cond_br24_falseOut_ready
    );

  cond_br25 : entity work.cond_br_dataless(arch)
    port map(
      condition => buffer134_outs,
      condition_valid => buffer134_outs_valid,
      condition_ready => buffer134_outs_ready,
      data_valid => cond_br22_falseOut_valid,
      data_ready => cond_br22_falseOut_ready,
      clk => clk,
      rst => rst,
      trueOut_valid => cond_br25_trueOut_valid,
      trueOut_ready => cond_br25_trueOut_ready,
      falseOut_valid => cond_br25_falseOut_valid,
      falseOut_ready => cond_br25_falseOut_ready
    );

  buffer134 : entity work.tfifo(arch) generic map(1, 1)
    port map(
      ins => fork53_outs_5,
      ins_valid => fork53_outs_5_valid,
      ins_ready => fork53_outs_5_ready,
      clk => clk,
      rst => rst,
      outs => buffer134_outs,
      outs_valid => buffer134_outs_valid,
      outs_ready => buffer134_outs_ready
    );

  cond_br126 : entity work.cond_br_dataless(arch)
    port map(
      condition => fork56_outs_2,
      condition_valid => fork56_outs_2_valid,
      condition_ready => fork56_outs_2_ready,
      data_valid => cond_br124_falseOut_valid,
      data_ready => cond_br124_falseOut_ready,
      clk => clk,
      rst => rst,
      trueOut_valid => cond_br126_trueOut_valid,
      trueOut_ready => cond_br126_trueOut_ready,
      falseOut_valid => cond_br126_falseOut_valid,
      falseOut_ready => cond_br126_falseOut_ready
    );

  sink14 : entity work.sink_dataless(arch)
    port map(
      ins_valid => cond_br126_trueOut_valid,
      ins_ready => cond_br126_trueOut_ready,
      clk => clk,
      rst => rst
    );

  cond_br127 : entity work.cond_br_dataless(arch)
    port map(
      condition => buffer136_outs,
      condition_valid => buffer136_outs_valid,
      condition_ready => buffer136_outs_ready,
      data_valid => cond_br125_falseOut_valid,
      data_ready => cond_br125_falseOut_ready,
      clk => clk,
      rst => rst,
      trueOut_valid => cond_br127_trueOut_valid,
      trueOut_ready => cond_br127_trueOut_ready,
      falseOut_valid => cond_br127_falseOut_valid,
      falseOut_ready => cond_br127_falseOut_ready
    );

  buffer136 : entity work.tfifo(arch) generic map(1, 1)
    port map(
      ins => fork56_outs_1,
      ins_valid => fork56_outs_1_valid,
      ins_ready => fork56_outs_1_ready,
      clk => clk,
      rst => rst,
      outs => buffer136_outs,
      outs_valid => buffer136_outs_valid,
      outs_ready => buffer136_outs_ready
    );

  buffer135 : entity work.oehb(arch) generic map(5)
    port map(
      ins => cond_br24_falseOut,
      ins_valid => cond_br24_falseOut_valid,
      ins_ready => cond_br24_falseOut_ready,
      clk => clk,
      rst => rst,
      outs => buffer135_outs,
      outs_valid => buffer135_outs_valid,
      outs_ready => buffer135_outs_ready
    );

  extsi83 : entity work.extsi(arch) generic map(5, 6)
    port map(
      ins => buffer135_outs,
      ins_valid => buffer135_outs_valid,
      ins_ready => buffer135_outs_ready,
      clk => clk,
      rst => rst,
      outs => extsi83_outs,
      outs_valid => extsi83_outs_valid,
      outs_ready => extsi83_outs_ready
    );

  fork54 : entity work.fork_dataless(arch) generic map(2)
    port map(
      ins_valid => cond_br25_falseOut_valid,
      ins_ready => cond_br25_falseOut_ready,
      clk => clk,
      rst => rst,
      outs_valid(0) => fork54_outs_0_valid,
      outs_valid(1) => fork54_outs_1_valid,
      outs_ready(0) => fork54_outs_0_ready,
      outs_ready(1) => fork54_outs_1_ready
    );

  constant71 : entity work.handshake_constant_0(arch) generic map(1)
    port map(
      ctrl_valid => fork54_outs_0_valid,
      ctrl_ready => fork54_outs_0_ready,
      clk => clk,
      rst => rst,
      outs => constant71_outs,
      outs_valid => constant71_outs_valid,
      outs_ready => constant71_outs_ready
    );

  source16 : entity work.source(arch)
    port map(
      clk => clk,
      rst => rst,
      outs_valid => source16_outs_valid,
      outs_ready => source16_outs_ready
    );

  constant72 : entity work.handshake_constant_3(arch) generic map(5)
    port map(
      ctrl_valid => source16_outs_valid,
      ctrl_ready => source16_outs_ready,
      clk => clk,
      rst => rst,
      outs => constant72_outs,
      outs_valid => constant72_outs_valid,
      outs_ready => constant72_outs_ready
    );

  extsi84 : entity work.extsi(arch) generic map(5, 6)
    port map(
      ins => constant72_outs,
      ins_valid => constant72_outs_valid,
      ins_ready => constant72_outs_ready,
      clk => clk,
      rst => rst,
      outs => extsi84_outs,
      outs_valid => extsi84_outs_valid,
      outs_ready => extsi84_outs_ready
    );

  source17 : entity work.source(arch)
    port map(
      clk => clk,
      rst => rst,
      outs_valid => source17_outs_valid,
      outs_ready => source17_outs_ready
    );

  constant73 : entity work.handshake_constant_1(arch) generic map(2)
    port map(
      ctrl_valid => source17_outs_valid,
      ctrl_ready => source17_outs_ready,
      clk => clk,
      rst => rst,
      outs => constant73_outs,
      outs_valid => constant73_outs_valid,
      outs_ready => constant73_outs_ready
    );

  extsi85 : entity work.extsi(arch) generic map(2, 6)
    port map(
      ins => constant73_outs,
      ins_valid => constant73_outs_valid,
      ins_ready => constant73_outs_ready,
      clk => clk,
      rst => rst,
      outs => extsi85_outs,
      outs_valid => extsi85_outs_valid,
      outs_ready => extsi85_outs_ready
    );

  addi23 : entity work.addi(arch) generic map(6)
    port map(
      lhs => extsi83_outs,
      lhs_valid => extsi83_outs_valid,
      lhs_ready => extsi83_outs_ready,
      rhs => extsi85_outs,
      rhs_valid => extsi85_outs_valid,
      rhs_ready => extsi85_outs_ready,
      clk => clk,
      rst => rst,
      result => addi23_result,
      result_valid => addi23_result_valid,
      result_ready => addi23_result_ready
    );

  buffer137 : entity work.oehb(arch) generic map(6)
    port map(
      ins => addi23_result,
      ins_valid => addi23_result_valid,
      ins_ready => addi23_result_ready,
      clk => clk,
      rst => rst,
      outs => buffer137_outs,
      outs_valid => buffer137_outs_valid,
      outs_ready => buffer137_outs_ready
    );

  fork55 : entity work.handshake_fork(arch) generic map(2, 6)
    port map(
      ins => buffer137_outs,
      ins_valid => buffer137_outs_valid,
      ins_ready => buffer137_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork55_outs_0,
      outs(1) => fork55_outs_1,
      outs_valid(0) => fork55_outs_0_valid,
      outs_valid(1) => fork55_outs_1_valid,
      outs_ready(0) => fork55_outs_0_ready,
      outs_ready(1) => fork55_outs_1_ready
    );

  trunci21 : entity work.trunci(arch) generic map(6, 5)
    port map(
      ins => fork55_outs_0,
      ins_valid => fork55_outs_0_valid,
      ins_ready => fork55_outs_0_ready,
      clk => clk,
      rst => rst,
      outs => trunci21_outs,
      outs_valid => trunci21_outs_valid,
      outs_ready => trunci21_outs_ready
    );

  cmpi5 : entity work.handshake_cmpi_0(arch) generic map(6)
    port map(
      lhs => fork55_outs_1,
      lhs_valid => fork55_outs_1_valid,
      lhs_ready => fork55_outs_1_ready,
      rhs => extsi84_outs,
      rhs_valid => extsi84_outs_valid,
      rhs_ready => extsi84_outs_ready,
      clk => clk,
      rst => rst,
      result => cmpi5_result,
      result_valid => cmpi5_result_valid,
      result_ready => cmpi5_result_ready
    );

  buffer138 : entity work.oehb(arch) generic map(1)
    port map(
      ins => cmpi5_result,
      ins_valid => cmpi5_result_valid,
      ins_ready => cmpi5_result_ready,
      clk => clk,
      rst => rst,
      outs => buffer138_outs,
      outs_valid => buffer138_outs_valid,
      outs_ready => buffer138_outs_ready
    );

  fork56 : entity work.handshake_fork(arch) generic map(6, 1)
    port map(
      ins => buffer138_outs,
      ins_valid => buffer138_outs_valid,
      ins_ready => buffer138_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork56_outs_0,
      outs(1) => fork56_outs_1,
      outs(2) => fork56_outs_2,
      outs(3) => fork56_outs_3,
      outs(4) => fork56_outs_4,
      outs(5) => fork56_outs_5,
      outs_valid(0) => fork56_outs_0_valid,
      outs_valid(1) => fork56_outs_1_valid,
      outs_valid(2) => fork56_outs_2_valid,
      outs_valid(3) => fork56_outs_3_valid,
      outs_valid(4) => fork56_outs_4_valid,
      outs_valid(5) => fork56_outs_5_valid,
      outs_ready(0) => fork56_outs_0_ready,
      outs_ready(1) => fork56_outs_1_ready,
      outs_ready(2) => fork56_outs_2_ready,
      outs_ready(3) => fork56_outs_3_ready,
      outs_ready(4) => fork56_outs_4_ready,
      outs_ready(5) => fork56_outs_5_ready
    );

  cond_br26 : entity work.cond_br(arch) generic map(5)
    port map(
      condition => fork56_outs_0,
      condition_valid => fork56_outs_0_valid,
      condition_ready => fork56_outs_0_ready,
      data => trunci21_outs,
      data_valid => trunci21_outs_valid,
      data_ready => trunci21_outs_ready,
      clk => clk,
      rst => rst,
      trueOut => cond_br26_trueOut,
      trueOut_valid => cond_br26_trueOut_valid,
      trueOut_ready => cond_br26_trueOut_ready,
      falseOut => cond_br26_falseOut,
      falseOut_valid => cond_br26_falseOut_valid,
      falseOut_ready => cond_br26_falseOut_ready
    );

  sink16 : entity work.sink(arch) generic map(5)
    port map(
      ins => cond_br26_falseOut,
      ins_valid => cond_br26_falseOut_valid,
      ins_ready => cond_br26_falseOut_ready,
      clk => clk,
      rst => rst
    );

  cond_br27 : entity work.cond_br_dataless(arch)
    port map(
      condition => fork56_outs_4,
      condition_valid => fork56_outs_4_valid,
      condition_ready => fork56_outs_4_ready,
      data_valid => fork54_outs_1_valid,
      data_ready => fork54_outs_1_ready,
      clk => clk,
      rst => rst,
      trueOut_valid => cond_br27_trueOut_valid,
      trueOut_ready => cond_br27_trueOut_ready,
      falseOut_valid => cond_br27_falseOut_valid,
      falseOut_ready => cond_br27_falseOut_ready
    );

  cond_br28 : entity work.cond_br(arch) generic map(1)
    port map(
      condition => fork56_outs_5,
      condition_valid => fork56_outs_5_valid,
      condition_ready => fork56_outs_5_ready,
      data => constant71_outs,
      data_valid => constant71_outs_valid,
      data_ready => constant71_outs_ready,
      clk => clk,
      rst => rst,
      trueOut => cond_br28_trueOut,
      trueOut_valid => cond_br28_trueOut_valid,
      trueOut_ready => cond_br28_trueOut_ready,
      falseOut => cond_br28_falseOut,
      falseOut_valid => cond_br28_falseOut_valid,
      falseOut_ready => cond_br28_falseOut_ready
    );

  sink17 : entity work.sink(arch) generic map(1)
    port map(
      ins => cond_br28_trueOut,
      ins_valid => cond_br28_trueOut_valid,
      ins_ready => cond_br28_trueOut_ready,
      clk => clk,
      rst => rst
    );

  extsi47 : entity work.extsi(arch) generic map(1, 5)
    port map(
      ins => cond_br28_falseOut,
      ins_valid => cond_br28_falseOut_valid,
      ins_ready => cond_br28_falseOut_ready,
      clk => clk,
      rst => rst,
      outs => extsi47_outs,
      outs_valid => extsi47_outs_valid,
      outs_ready => extsi47_outs_ready
    );

  init28 : entity work.tehb_init(arch) generic map(1, 0)
    port map(
      ins => fork96_outs_6,
      ins_valid => fork96_outs_6_valid,
      ins_ready => fork96_outs_6_ready,
      clk => clk,
      rst => rst,
      outs => init28_outs,
      outs_valid => init28_outs_valid,
      outs_ready => init28_outs_ready
    );

  fork57 : entity work.handshake_fork(arch) generic map(5, 1)
    port map(
      ins => init28_outs,
      ins_valid => init28_outs_valid,
      ins_ready => init28_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork57_outs_0,
      outs(1) => fork57_outs_1,
      outs(2) => fork57_outs_2,
      outs(3) => fork57_outs_3,
      outs(4) => fork57_outs_4,
      outs_valid(0) => fork57_outs_0_valid,
      outs_valid(1) => fork57_outs_1_valid,
      outs_valid(2) => fork57_outs_2_valid,
      outs_valid(3) => fork57_outs_3_valid,
      outs_valid(4) => fork57_outs_4_valid,
      outs_ready(0) => fork57_outs_0_ready,
      outs_ready(1) => fork57_outs_1_ready,
      outs_ready(2) => fork57_outs_2_ready,
      outs_ready(3) => fork57_outs_3_ready,
      outs_ready(4) => fork57_outs_4_ready
    );

  mux46 : entity work.mux_dataless(arch) generic map(2, 1)
    port map(
      index => buffer143_outs,
      index_valid => buffer143_outs_valid,
      index_ready => buffer143_outs_ready,
      ins_valid(0) => cond_br126_falseOut_valid,
      ins_valid(1) => cond_br139_trueOut_valid,
      ins_ready(0) => cond_br126_falseOut_ready,
      ins_ready(1) => cond_br139_trueOut_ready,
      clk => clk,
      rst => rst,
      outs_valid => mux46_outs_valid,
      outs_ready => mux46_outs_ready
    );

  buffer143 : entity work.tfifo(arch) generic map(1, 1)
    port map(
      ins => fork57_outs_4,
      ins_valid => fork57_outs_4_valid,
      ins_ready => fork57_outs_4_ready,
      clk => clk,
      rst => rst,
      outs => buffer143_outs,
      outs_valid => buffer143_outs_valid,
      outs_ready => buffer143_outs_ready
    );

  buffer139 : entity work.oehb_dataless(arch)
    port map(
      ins_valid => mux46_outs_valid,
      ins_ready => mux46_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer139_outs_valid,
      outs_ready => buffer139_outs_ready
    );

  buffer140 : entity work.tehb_dataless(arch)
    port map(
      ins_valid => buffer139_outs_valid,
      ins_ready => buffer139_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer140_outs_valid,
      outs_ready => buffer140_outs_ready
    );

  fork58 : entity work.fork_dataless(arch) generic map(2)
    port map(
      ins_valid => buffer140_outs_valid,
      ins_ready => buffer140_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid(0) => fork58_outs_0_valid,
      outs_valid(1) => fork58_outs_1_valid,
      outs_ready(0) => fork58_outs_0_ready,
      outs_ready(1) => fork58_outs_1_ready
    );

  mux47 : entity work.mux_dataless(arch) generic map(2, 1)
    port map(
      index => buffer144_outs,
      index_valid => buffer144_outs_valid,
      index_ready => buffer144_outs_ready,
      ins_valid(0) => cond_br127_falseOut_valid,
      ins_valid(1) => cond_br142_trueOut_valid,
      ins_ready(0) => cond_br127_falseOut_ready,
      ins_ready(1) => cond_br142_trueOut_ready,
      clk => clk,
      rst => rst,
      outs_valid => mux47_outs_valid,
      outs_ready => mux47_outs_ready
    );

  buffer144 : entity work.tfifo(arch) generic map(1, 1)
    port map(
      ins => fork57_outs_3,
      ins_valid => fork57_outs_3_valid,
      ins_ready => fork57_outs_3_ready,
      clk => clk,
      rst => rst,
      outs => buffer144_outs,
      outs_valid => buffer144_outs_valid,
      outs_ready => buffer144_outs_ready
    );

  buffer141 : entity work.oehb_dataless(arch)
    port map(
      ins_valid => mux47_outs_valid,
      ins_ready => mux47_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer141_outs_valid,
      outs_ready => buffer141_outs_ready
    );

  buffer142 : entity work.tehb_dataless(arch)
    port map(
      ins_valid => buffer141_outs_valid,
      ins_ready => buffer141_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer142_outs_valid,
      outs_ready => buffer142_outs_ready
    );

  fork59 : entity work.fork_dataless(arch) generic map(2)
    port map(
      ins_valid => buffer142_outs_valid,
      ins_ready => buffer142_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid(0) => fork59_outs_0_valid,
      outs_valid(1) => fork59_outs_1_valid,
      outs_ready(0) => fork59_outs_0_ready,
      outs_ready(1) => fork59_outs_1_ready
    );

  buffer245 : entity work.oehb_dataless(arch)
    port map(
      ins_valid => cond_br141_trueOut_valid,
      ins_ready => cond_br141_trueOut_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer245_outs_valid,
      outs_ready => buffer245_outs_ready
    );

  mux48 : entity work.mux_dataless(arch) generic map(2, 1)
    port map(
      index => buffer145_outs,
      index_valid => buffer145_outs_valid,
      index_ready => buffer145_outs_ready,
      ins_valid(0) => cond_br120_falseOut_valid,
      ins_valid(1) => buffer245_outs_valid,
      ins_ready(0) => cond_br120_falseOut_ready,
      ins_ready(1) => buffer245_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => mux48_outs_valid,
      outs_ready => mux48_outs_ready
    );

  buffer145 : entity work.tfifo(arch) generic map(1, 1)
    port map(
      ins => fork57_outs_2,
      ins_valid => fork57_outs_2_valid,
      ins_ready => fork57_outs_2_ready,
      clk => clk,
      rst => rst,
      outs => buffer145_outs,
      outs_valid => buffer145_outs_valid,
      outs_ready => buffer145_outs_ready
    );

  buffer146 : entity work.tehb_dataless(arch)
    port map(
      ins_valid => mux48_outs_valid,
      ins_ready => mux48_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer146_outs_valid,
      outs_ready => buffer146_outs_ready
    );

  fork60 : entity work.fork_dataless(arch) generic map(2)
    port map(
      ins_valid => buffer146_outs_valid,
      ins_ready => buffer146_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid(0) => fork60_outs_0_valid,
      outs_valid(1) => fork60_outs_1_valid,
      outs_ready(0) => fork60_outs_0_ready,
      outs_ready(1) => fork60_outs_1_ready
    );

  mux49 : entity work.mux_dataless(arch) generic map(2, 1)
    port map(
      index => fork57_outs_1,
      index_valid => fork57_outs_1_valid,
      index_ready => fork57_outs_1_ready,
      ins_valid(0) => cond_br121_falseOut_valid,
      ins_valid(1) => cond_br143_trueOut_valid,
      ins_ready(0) => cond_br121_falseOut_ready,
      ins_ready(1) => cond_br143_trueOut_ready,
      clk => clk,
      rst => rst,
      outs_valid => mux49_outs_valid,
      outs_ready => mux49_outs_ready
    );

  buffer147 : entity work.oehb_dataless(arch)
    port map(
      ins_valid => mux49_outs_valid,
      ins_ready => mux49_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer147_outs_valid,
      outs_ready => buffer147_outs_ready
    );

  buffer148 : entity work.tehb_dataless(arch)
    port map(
      ins_valid => buffer147_outs_valid,
      ins_ready => buffer147_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer148_outs_valid,
      outs_ready => buffer148_outs_ready
    );

  fork61 : entity work.fork_dataless(arch) generic map(2)
    port map(
      ins_valid => buffer148_outs_valid,
      ins_ready => buffer148_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid(0) => fork61_outs_0_valid,
      outs_valid(1) => fork61_outs_1_valid,
      outs_ready(0) => fork61_outs_0_ready,
      outs_ready(1) => fork61_outs_1_ready
    );

  mux51 : entity work.mux_dataless(arch) generic map(2, 1)
    port map(
      index => fork57_outs_0,
      index_valid => fork57_outs_0_valid,
      index_ready => fork57_outs_0_ready,
      ins_valid(0) => fork0_outs_2_valid,
      ins_valid(1) => cond_br140_trueOut_valid,
      ins_ready(0) => fork0_outs_2_ready,
      ins_ready(1) => cond_br140_trueOut_ready,
      clk => clk,
      rst => rst,
      outs_valid => mux51_outs_valid,
      outs_ready => mux51_outs_ready
    );

  mux12 : entity work.mux(arch) generic map(2, 5, 1)
    port map(
      index => control_merge10_index,
      index_valid => control_merge10_index_valid,
      index_ready => control_merge10_index_ready,
      ins(0) => extsi47_outs,
      ins(1) => cond_br36_trueOut,
      ins_valid(0) => extsi47_outs_valid,
      ins_valid(1) => cond_br36_trueOut_valid,
      ins_ready(0) => extsi47_outs_ready,
      ins_ready(1) => cond_br36_trueOut_ready,
      clk => clk,
      rst => rst,
      outs => mux12_outs,
      outs_valid => mux12_outs_valid,
      outs_ready => mux12_outs_ready
    );

  control_merge10 : entity work.control_merge_dataless(arch) generic map(2, 1)
    port map(
      ins_valid(0) => cond_br27_falseOut_valid,
      ins_valid(1) => cond_br37_trueOut_valid,
      ins_ready(0) => cond_br27_falseOut_ready,
      ins_ready(1) => cond_br37_trueOut_ready,
      clk => clk,
      rst => rst,
      outs_valid => control_merge10_outs_valid,
      outs_ready => control_merge10_outs_ready,
      index => control_merge10_index,
      index_valid => control_merge10_index_valid,
      index_ready => control_merge10_index_ready
    );

  fork62 : entity work.fork_dataless(arch) generic map(2)
    port map(
      ins_valid => control_merge10_outs_valid,
      ins_ready => control_merge10_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid(0) => fork62_outs_0_valid,
      outs_valid(1) => fork62_outs_1_valid,
      outs_ready(0) => fork62_outs_0_ready,
      outs_ready(1) => fork62_outs_1_ready
    );

  constant74 : entity work.handshake_constant_0(arch) generic map(1)
    port map(
      ctrl_valid => fork62_outs_0_valid,
      ctrl_ready => fork62_outs_0_ready,
      clk => clk,
      rst => rst,
      outs => constant74_outs,
      outs_valid => constant74_outs_valid,
      outs_ready => constant74_outs_ready
    );

  extsi46 : entity work.extsi(arch) generic map(1, 5)
    port map(
      ins => constant74_outs,
      ins_valid => constant74_outs_valid,
      ins_ready => constant74_outs_ready,
      clk => clk,
      rst => rst,
      outs => extsi46_outs,
      outs_valid => extsi46_outs_valid,
      outs_ready => extsi46_outs_ready
    );

  buffer151 : entity work.tehb(arch) generic map(5)
    port map(
      ins => mux12_outs,
      ins_valid => mux12_outs_valid,
      ins_ready => mux12_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer151_outs,
      outs_valid => buffer151_outs_valid,
      outs_ready => buffer151_outs_ready
    );

  init35 : entity work.tehb_init(arch) generic map(1, 0)
    port map(
      ins => fork94_outs_7,
      ins_valid => fork94_outs_7_valid,
      ins_ready => fork94_outs_7_ready,
      clk => clk,
      rst => rst,
      outs => init35_outs,
      outs_valid => init35_outs_valid,
      outs_ready => init35_outs_ready
    );

  fork63 : entity work.handshake_fork(arch) generic map(5, 1)
    port map(
      ins => init35_outs,
      ins_valid => init35_outs_valid,
      ins_ready => init35_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork63_outs_0,
      outs(1) => fork63_outs_1,
      outs(2) => fork63_outs_2,
      outs(3) => fork63_outs_3,
      outs(4) => fork63_outs_4,
      outs_valid(0) => fork63_outs_0_valid,
      outs_valid(1) => fork63_outs_1_valid,
      outs_valid(2) => fork63_outs_2_valid,
      outs_valid(3) => fork63_outs_3_valid,
      outs_valid(4) => fork63_outs_4_valid,
      outs_ready(0) => fork63_outs_0_ready,
      outs_ready(1) => fork63_outs_1_ready,
      outs_ready(2) => fork63_outs_2_ready,
      outs_ready(3) => fork63_outs_3_ready,
      outs_ready(4) => fork63_outs_4_ready
    );

  mux53 : entity work.mux_dataless(arch) generic map(2, 1)
    port map(
      index => fork63_outs_4,
      index_valid => fork63_outs_4_valid,
      index_ready => fork63_outs_4_ready,
      ins_valid(0) => fork58_outs_1_valid,
      ins_valid(1) => cond_br135_trueOut_valid,
      ins_ready(0) => fork58_outs_1_ready,
      ins_ready(1) => cond_br135_trueOut_ready,
      clk => clk,
      rst => rst,
      outs_valid => mux53_outs_valid,
      outs_ready => mux53_outs_ready
    );

  buffer152 : entity work.oehb_dataless(arch)
    port map(
      ins_valid => mux53_outs_valid,
      ins_ready => mux53_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer152_outs_valid,
      outs_ready => buffer152_outs_ready
    );

  buffer154 : entity work.tehb_dataless(arch)
    port map(
      ins_valid => buffer152_outs_valid,
      ins_ready => buffer152_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer154_outs_valid,
      outs_ready => buffer154_outs_ready
    );

  fork64 : entity work.fork_dataless(arch) generic map(2)
    port map(
      ins_valid => buffer154_outs_valid,
      ins_ready => buffer154_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid(0) => fork64_outs_0_valid,
      outs_valid(1) => fork64_outs_1_valid,
      outs_ready(0) => fork64_outs_0_ready,
      outs_ready(1) => fork64_outs_1_ready
    );

  buffer242 : entity work.oehb_dataless(arch)
    port map(
      ins_valid => cond_br137_trueOut_valid,
      ins_ready => cond_br137_trueOut_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer242_outs_valid,
      outs_ready => buffer242_outs_ready
    );

  mux54 : entity work.mux_dataless(arch) generic map(2, 1)
    port map(
      index => fork63_outs_3,
      index_valid => fork63_outs_3_valid,
      index_ready => fork63_outs_3_ready,
      ins_valid(0) => fork59_outs_1_valid,
      ins_valid(1) => buffer242_outs_valid,
      ins_ready(0) => fork59_outs_1_ready,
      ins_ready(1) => buffer242_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => mux54_outs_valid,
      outs_ready => mux54_outs_ready
    );

  buffer155 : entity work.tehb_dataless(arch)
    port map(
      ins_valid => mux54_outs_valid,
      ins_ready => mux54_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer155_outs_valid,
      outs_ready => buffer155_outs_ready
    );

  fork65 : entity work.fork_dataless(arch) generic map(2)
    port map(
      ins_valid => buffer155_outs_valid,
      ins_ready => buffer155_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid(0) => fork65_outs_0_valid,
      outs_valid(1) => fork65_outs_1_valid,
      outs_ready(0) => fork65_outs_0_ready,
      outs_ready(1) => fork65_outs_1_ready
    );

  mux55 : entity work.mux_dataless(arch) generic map(2, 1)
    port map(
      index => fork63_outs_2,
      index_valid => fork63_outs_2_valid,
      index_ready => fork63_outs_2_ready,
      ins_valid(0) => fork60_outs_1_valid,
      ins_valid(1) => cond_br138_trueOut_valid,
      ins_ready(0) => fork60_outs_1_ready,
      ins_ready(1) => cond_br138_trueOut_ready,
      clk => clk,
      rst => rst,
      outs_valid => mux55_outs_valid,
      outs_ready => mux55_outs_ready
    );

  buffer156 : entity work.oehb_dataless(arch)
    port map(
      ins_valid => mux55_outs_valid,
      ins_ready => mux55_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer156_outs_valid,
      outs_ready => buffer156_outs_ready
    );

  buffer157 : entity work.tehb_dataless(arch)
    port map(
      ins_valid => buffer156_outs_valid,
      ins_ready => buffer156_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer157_outs_valid,
      outs_ready => buffer157_outs_ready
    );

  fork66 : entity work.fork_dataless(arch) generic map(2)
    port map(
      ins_valid => buffer157_outs_valid,
      ins_ready => buffer157_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid(0) => fork66_outs_0_valid,
      outs_valid(1) => fork66_outs_1_valid,
      outs_ready(0) => fork66_outs_0_ready,
      outs_ready(1) => fork66_outs_1_ready
    );

  mux56 : entity work.mux_dataless(arch) generic map(2, 1)
    port map(
      index => fork63_outs_1,
      index_valid => fork63_outs_1_valid,
      index_ready => fork63_outs_1_ready,
      ins_valid(0) => fork61_outs_1_valid,
      ins_valid(1) => cond_br136_trueOut_valid,
      ins_ready(0) => fork61_outs_1_ready,
      ins_ready(1) => cond_br136_trueOut_ready,
      clk => clk,
      rst => rst,
      outs_valid => mux56_outs_valid,
      outs_ready => mux56_outs_ready
    );

  buffer158 : entity work.oehb_dataless(arch)
    port map(
      ins_valid => mux56_outs_valid,
      ins_ready => mux56_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer158_outs_valid,
      outs_ready => buffer158_outs_ready
    );

  buffer159 : entity work.tehb_dataless(arch)
    port map(
      ins_valid => buffer158_outs_valid,
      ins_ready => buffer158_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer159_outs_valid,
      outs_ready => buffer159_outs_ready
    );

  fork67 : entity work.fork_dataless(arch) generic map(2)
    port map(
      ins_valid => buffer159_outs_valid,
      ins_ready => buffer159_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid(0) => fork67_outs_0_valid,
      outs_valid(1) => fork67_outs_1_valid,
      outs_ready(0) => fork67_outs_0_ready,
      outs_ready(1) => fork67_outs_1_ready
    );

  buffer149 : entity work.oehb_dataless(arch)
    port map(
      ins_valid => mux51_outs_valid,
      ins_ready => mux51_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer149_outs_valid,
      outs_ready => buffer149_outs_ready
    );

  buffer150 : entity work.tehb_dataless(arch)
    port map(
      ins_valid => buffer149_outs_valid,
      ins_ready => buffer149_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer150_outs_valid,
      outs_ready => buffer150_outs_ready
    );

  mux58 : entity work.mux_dataless(arch) generic map(2, 1)
    port map(
      index => buffer153_outs,
      index_valid => buffer153_outs_valid,
      index_ready => buffer153_outs_ready,
      ins_valid(0) => buffer150_outs_valid,
      ins_valid(1) => cond_br134_trueOut_valid,
      ins_ready(0) => buffer150_outs_ready,
      ins_ready(1) => cond_br134_trueOut_ready,
      clk => clk,
      rst => rst,
      outs_valid => mux58_outs_valid,
      outs_ready => mux58_outs_ready
    );

  buffer153 : entity work.tfifo(arch) generic map(1, 1)
    port map(
      ins => fork63_outs_0,
      ins_valid => fork63_outs_0_valid,
      ins_ready => fork63_outs_0_ready,
      clk => clk,
      rst => rst,
      outs => buffer153_outs,
      outs_valid => buffer153_outs_valid,
      outs_ready => buffer153_outs_ready
    );

  mux13 : entity work.mux(arch) generic map(2, 5, 1)
    port map(
      index => fork71_outs_1,
      index_valid => fork71_outs_1_valid,
      index_ready => fork71_outs_1_ready,
      ins(0) => extsi46_outs,
      ins(1) => cond_br33_trueOut,
      ins_valid(0) => extsi46_outs_valid,
      ins_valid(1) => cond_br33_trueOut_valid,
      ins_ready(0) => extsi46_outs_ready,
      ins_ready(1) => cond_br33_trueOut_ready,
      clk => clk,
      rst => rst,
      outs => mux13_outs,
      outs_valid => mux13_outs_valid,
      outs_ready => mux13_outs_ready
    );

  buffer161 : entity work.tehb(arch) generic map(5)
    port map(
      ins => mux13_outs,
      ins_valid => mux13_outs_valid,
      ins_ready => mux13_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer161_outs,
      outs_valid => buffer161_outs_valid,
      outs_ready => buffer161_outs_ready
    );

  fork68 : entity work.handshake_fork(arch) generic map(2, 5)
    port map(
      ins => buffer161_outs,
      ins_valid => buffer161_outs_valid,
      ins_ready => buffer161_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork68_outs_0,
      outs(1) => fork68_outs_1,
      outs_valid(0) => fork68_outs_0_valid,
      outs_valid(1) => fork68_outs_1_valid,
      outs_ready(0) => fork68_outs_0_ready,
      outs_ready(1) => fork68_outs_1_ready
    );

  extsi86 : entity work.extsi(arch) generic map(5, 7)
    port map(
      ins => fork68_outs_0,
      ins_valid => fork68_outs_0_valid,
      ins_ready => fork68_outs_0_ready,
      clk => clk,
      rst => rst,
      outs => extsi86_outs,
      outs_valid => extsi86_outs_valid,
      outs_ready => extsi86_outs_ready
    );

  mux14 : entity work.mux(arch) generic map(2, 5, 1)
    port map(
      index => fork71_outs_0,
      index_valid => fork71_outs_0_valid,
      index_ready => fork71_outs_0_ready,
      ins(0) => buffer151_outs,
      ins(1) => cond_br34_trueOut,
      ins_valid(0) => buffer151_outs_valid,
      ins_valid(1) => cond_br34_trueOut_valid,
      ins_ready(0) => buffer151_outs_ready,
      ins_ready(1) => cond_br34_trueOut_ready,
      clk => clk,
      rst => rst,
      outs => mux14_outs,
      outs_valid => mux14_outs_valid,
      outs_ready => mux14_outs_ready
    );

  buffer162 : entity work.oehb(arch) generic map(5)
    port map(
      ins => mux14_outs,
      ins_valid => mux14_outs_valid,
      ins_ready => mux14_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer162_outs,
      outs_valid => buffer162_outs_valid,
      outs_ready => buffer162_outs_ready
    );

  buffer163 : entity work.tehb(arch) generic map(5)
    port map(
      ins => buffer162_outs,
      ins_valid => buffer162_outs_valid,
      ins_ready => buffer162_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer163_outs,
      outs_valid => buffer163_outs_valid,
      outs_ready => buffer163_outs_ready
    );

  fork69 : entity work.handshake_fork(arch) generic map(2, 5)
    port map(
      ins => buffer163_outs,
      ins_valid => buffer163_outs_valid,
      ins_ready => buffer163_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork69_outs_0,
      outs(1) => fork69_outs_1,
      outs_valid(0) => fork69_outs_0_valid,
      outs_valid(1) => fork69_outs_1_valid,
      outs_ready(0) => fork69_outs_0_ready,
      outs_ready(1) => fork69_outs_1_ready
    );

  extsi87 : entity work.extsi(arch) generic map(5, 32)
    port map(
      ins => fork69_outs_1,
      ins_valid => fork69_outs_1_valid,
      ins_ready => fork69_outs_1_ready,
      clk => clk,
      rst => rst,
      outs => extsi87_outs,
      outs_valid => extsi87_outs_valid,
      outs_ready => extsi87_outs_ready
    );

  fork70 : entity work.handshake_fork(arch) generic map(2, 32)
    port map(
      ins => extsi87_outs,
      ins_valid => extsi87_outs_valid,
      ins_ready => extsi87_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork70_outs_0,
      outs(1) => fork70_outs_1,
      outs_valid(0) => fork70_outs_0_valid,
      outs_valid(1) => fork70_outs_1_valid,
      outs_ready(0) => fork70_outs_0_ready,
      outs_ready(1) => fork70_outs_1_ready
    );

  control_merge11 : entity work.control_merge_dataless(arch) generic map(2, 1)
    port map(
      ins_valid(0) => fork62_outs_1_valid,
      ins_valid(1) => cond_br35_trueOut_valid,
      ins_ready(0) => fork62_outs_1_ready,
      ins_ready(1) => cond_br35_trueOut_ready,
      clk => clk,
      rst => rst,
      outs_valid => control_merge11_outs_valid,
      outs_ready => control_merge11_outs_ready,
      index => control_merge11_index,
      index_valid => control_merge11_index_valid,
      index_ready => control_merge11_index_ready
    );

  fork71 : entity work.handshake_fork(arch) generic map(2, 1)
    port map(
      ins => control_merge11_index,
      ins_valid => control_merge11_index_valid,
      ins_ready => control_merge11_index_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork71_outs_0,
      outs(1) => fork71_outs_1,
      outs_valid(0) => fork71_outs_0_valid,
      outs_valid(1) => fork71_outs_1_valid,
      outs_ready(0) => fork71_outs_0_ready,
      outs_ready(1) => fork71_outs_1_ready
    );

  fork72 : entity work.fork_dataless(arch) generic map(3)
    port map(
      ins_valid => control_merge11_outs_valid,
      ins_ready => control_merge11_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid(0) => fork72_outs_0_valid,
      outs_valid(1) => fork72_outs_1_valid,
      outs_valid(2) => fork72_outs_2_valid,
      outs_ready(0) => fork72_outs_0_ready,
      outs_ready(1) => fork72_outs_1_ready,
      outs_ready(2) => fork72_outs_2_ready
    );

  constant75 : entity work.handshake_constant_1(arch) generic map(2)
    port map(
      ctrl_valid => fork72_outs_1_valid,
      ctrl_ready => fork72_outs_1_ready,
      clk => clk,
      rst => rst,
      outs => constant75_outs,
      outs_valid => constant75_outs_valid,
      outs_ready => constant75_outs_ready
    );

  extsi32 : entity work.extsi(arch) generic map(2, 32)
    port map(
      ins => constant75_outs,
      ins_valid => constant75_outs_valid,
      ins_ready => constant75_outs_ready,
      clk => clk,
      rst => rst,
      outs => extsi32_outs,
      outs_valid => extsi32_outs_valid,
      outs_ready => extsi32_outs_ready
    );

  constant76 : entity work.handshake_constant_0(arch) generic map(1)
    port map(
      ctrl_valid => fork72_outs_0_valid,
      ctrl_ready => fork72_outs_0_ready,
      clk => clk,
      rst => rst,
      outs => constant76_outs,
      outs_valid => constant76_outs_valid,
      outs_ready => constant76_outs_ready
    );

  fork73 : entity work.handshake_fork(arch) generic map(2, 1)
    port map(
      ins => constant76_outs,
      ins_valid => constant76_outs_valid,
      ins_ready => constant76_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork73_outs_0,
      outs(1) => fork73_outs_1,
      outs_valid(0) => fork73_outs_0_valid,
      outs_valid(1) => fork73_outs_1_valid,
      outs_ready(0) => fork73_outs_0_ready,
      outs_ready(1) => fork73_outs_1_ready
    );

  extsi34 : entity work.extsi(arch) generic map(1, 32)
    port map(
      ins => fork73_outs_1,
      ins_valid => fork73_outs_1_valid,
      ins_ready => fork73_outs_1_ready,
      clk => clk,
      rst => rst,
      outs => extsi34_outs,
      outs_valid => extsi34_outs_valid,
      outs_ready => extsi34_outs_ready
    );

  source18 : entity work.source(arch)
    port map(
      clk => clk,
      rst => rst,
      outs_valid => source18_outs_valid,
      outs_ready => source18_outs_ready
    );

  constant77 : entity work.handshake_constant_1(arch) generic map(2)
    port map(
      ctrl_valid => source18_outs_valid,
      ctrl_ready => source18_outs_ready,
      clk => clk,
      rst => rst,
      outs => constant77_outs,
      outs_valid => constant77_outs_valid,
      outs_ready => constant77_outs_ready
    );

  extsi35 : entity work.extsi(arch) generic map(2, 32)
    port map(
      ins => constant77_outs,
      ins_valid => constant77_outs_valid,
      ins_ready => constant77_outs_ready,
      clk => clk,
      rst => rst,
      outs => extsi35_outs,
      outs_valid => extsi35_outs_valid,
      outs_ready => extsi35_outs_ready
    );

  source19 : entity work.source(arch)
    port map(
      clk => clk,
      rst => rst,
      outs_valid => source19_outs_valid,
      outs_ready => source19_outs_ready
    );

  constant78 : entity work.handshake_constant_2(arch) generic map(3)
    port map(
      ctrl_valid => source19_outs_valid,
      ctrl_ready => source19_outs_ready,
      clk => clk,
      rst => rst,
      outs => constant78_outs,
      outs_valid => constant78_outs_valid,
      outs_ready => constant78_outs_ready
    );

  extsi36 : entity work.extsi(arch) generic map(3, 32)
    port map(
      ins => constant78_outs,
      ins_valid => constant78_outs_valid,
      ins_ready => constant78_outs_ready,
      clk => clk,
      rst => rst,
      outs => extsi36_outs,
      outs_valid => extsi36_outs_valid,
      outs_ready => extsi36_outs_ready
    );

  shli20 : entity work.shli(arch) generic map(32)
    port map(
      lhs => fork70_outs_0,
      lhs_valid => fork70_outs_0_valid,
      lhs_ready => fork70_outs_0_ready,
      rhs => extsi35_outs,
      rhs_valid => extsi35_outs_valid,
      rhs_ready => extsi35_outs_ready,
      clk => clk,
      rst => rst,
      result => shli20_result,
      result_valid => shli20_result_valid,
      result_ready => shli20_result_ready
    );

  buffer170 : entity work.oehb(arch) generic map(32)
    port map(
      ins => shli20_result,
      ins_valid => shli20_result_valid,
      ins_ready => shli20_result_ready,
      clk => clk,
      rst => rst,
      outs => buffer170_outs,
      outs_valid => buffer170_outs_valid,
      outs_ready => buffer170_outs_ready
    );

  trunci22 : entity work.trunci(arch) generic map(32, 7)
    port map(
      ins => buffer170_outs,
      ins_valid => buffer170_outs_valid,
      ins_ready => buffer170_outs_ready,
      clk => clk,
      rst => rst,
      outs => trunci22_outs,
      outs_valid => trunci22_outs_valid,
      outs_ready => trunci22_outs_ready
    );

  shli21 : entity work.shli(arch) generic map(32)
    port map(
      lhs => fork70_outs_1,
      lhs_valid => fork70_outs_1_valid,
      lhs_ready => fork70_outs_1_ready,
      rhs => extsi36_outs,
      rhs_valid => extsi36_outs_valid,
      rhs_ready => extsi36_outs_ready,
      clk => clk,
      rst => rst,
      result => shli21_result,
      result_valid => shli21_result_valid,
      result_ready => shli21_result_ready
    );

  buffer177 : entity work.oehb(arch) generic map(32)
    port map(
      ins => shli21_result,
      ins_valid => shli21_result_valid,
      ins_ready => shli21_result_ready,
      clk => clk,
      rst => rst,
      outs => buffer177_outs,
      outs_valid => buffer177_outs_valid,
      outs_ready => buffer177_outs_ready
    );

  trunci23 : entity work.trunci(arch) generic map(32, 7)
    port map(
      ins => buffer177_outs,
      ins_valid => buffer177_outs_valid,
      ins_ready => buffer177_outs_ready,
      clk => clk,
      rst => rst,
      outs => trunci23_outs,
      outs_valid => trunci23_outs_valid,
      outs_ready => trunci23_outs_ready
    );

  addi37 : entity work.addi(arch) generic map(7)
    port map(
      lhs => trunci22_outs,
      lhs_valid => trunci22_outs_valid,
      lhs_ready => trunci22_outs_ready,
      rhs => trunci23_outs,
      rhs_valid => trunci23_outs_valid,
      rhs_ready => trunci23_outs_ready,
      clk => clk,
      rst => rst,
      result => addi37_result,
      result_valid => addi37_result_valid,
      result_ready => addi37_result_ready
    );

  buffer178 : entity work.oehb(arch) generic map(7)
    port map(
      ins => addi37_result,
      ins_valid => addi37_result_valid,
      ins_ready => addi37_result_ready,
      clk => clk,
      rst => rst,
      outs => buffer178_outs,
      outs_valid => buffer178_outs_valid,
      outs_ready => buffer178_outs_ready
    );

  addi13 : entity work.addi(arch) generic map(7)
    port map(
      lhs => extsi86_outs,
      lhs_valid => extsi86_outs_valid,
      lhs_ready => extsi86_outs_ready,
      rhs => buffer178_outs,
      rhs_valid => buffer178_outs_valid,
      rhs_ready => buffer178_outs_ready,
      clk => clk,
      rst => rst,
      result => addi13_result,
      result_valid => addi13_result_valid,
      result_ready => addi13_result_ready
    );

  buffer4 : entity work.tfifo_dataless(arch) generic map(1)
    port map(
      ins_valid => store4_doneOut_valid,
      ins_ready => store4_doneOut_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer4_outs_valid,
      outs_ready => buffer4_outs_ready
    );

  buffer179 : entity work.oehb(arch) generic map(7)
    port map(
      ins => addi13_result,
      ins_valid => addi13_result_valid,
      ins_ready => addi13_result_ready,
      clk => clk,
      rst => rst,
      outs => buffer179_outs,
      outs_valid => buffer179_outs_valid,
      outs_ready => buffer179_outs_ready
    );

  store4 : entity work.store(arch) generic map(32, 7)
    port map(
      addrIn => buffer179_outs,
      addrIn_valid => buffer179_outs_valid,
      addrIn_ready => buffer179_outs_ready,
      dataIn => extsi34_outs,
      dataIn_valid => extsi34_outs_valid,
      dataIn_ready => extsi34_outs_ready,
      doneFromMem_valid => mem_controller4_stDone_0_valid,
      doneFromMem_ready => mem_controller4_stDone_0_ready,
      clk => clk,
      rst => rst,
      addrOut => store4_addrOut,
      addrOut_valid => store4_addrOut_valid,
      addrOut_ready => store4_addrOut_ready,
      dataToMem => store4_dataToMem,
      dataToMem_valid => store4_dataToMem_valid,
      dataToMem_ready => store4_dataToMem_ready,
      doneOut_valid => store4_doneOut_valid,
      doneOut_ready => store4_doneOut_ready
    );

  extsi45 : entity work.extsi(arch) generic map(1, 5)
    port map(
      ins => fork73_outs_0,
      ins_valid => fork73_outs_0_valid,
      ins_ready => fork73_outs_0_ready,
      clk => clk,
      rst => rst,
      outs => extsi45_outs,
      outs_valid => extsi45_outs_valid,
      outs_ready => extsi45_outs_ready
    );

  buffer208 : entity work.oehb_dataless(arch)
    port map(
      ins_valid => fork79_outs_1_valid,
      ins_ready => fork79_outs_1_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer208_outs_valid,
      outs_ready => buffer208_outs_ready
    );

  cond_br128 : entity work.cond_br_dataless(arch)
    port map(
      condition => buffer164_outs,
      condition_valid => buffer164_outs_valid,
      condition_ready => buffer164_outs_ready,
      data_valid => buffer208_outs_valid,
      data_ready => buffer208_outs_ready,
      clk => clk,
      rst => rst,
      trueOut_valid => cond_br128_trueOut_valid,
      trueOut_ready => cond_br128_trueOut_ready,
      falseOut_valid => cond_br128_falseOut_valid,
      falseOut_ready => cond_br128_falseOut_ready
    );

  buffer164 : entity work.tfifo(arch) generic map(1, 1)
    port map(
      ins => fork92_outs_9,
      ins_valid => fork92_outs_9_valid,
      ins_ready => fork92_outs_9_ready,
      clk => clk,
      rst => rst,
      outs => buffer164_outs,
      outs_valid => buffer164_outs_valid,
      outs_ready => buffer164_outs_ready
    );

  sink18 : entity work.sink_dataless(arch)
    port map(
      ins_valid => cond_br128_falseOut_valid,
      ins_ready => cond_br128_falseOut_ready,
      clk => clk,
      rst => rst
    );

  cond_br129 : entity work.cond_br_dataless(arch)
    port map(
      condition => buffer165_outs,
      condition_valid => buffer165_outs_valid,
      condition_ready => buffer165_outs_ready,
      data_valid => fork75_outs_2_valid,
      data_ready => fork75_outs_2_ready,
      clk => clk,
      rst => rst,
      trueOut_valid => cond_br129_trueOut_valid,
      trueOut_ready => cond_br129_trueOut_ready,
      falseOut_valid => cond_br129_falseOut_valid,
      falseOut_ready => cond_br129_falseOut_ready
    );

  buffer165 : entity work.tfifo(arch) generic map(3, 1)
    port map(
      ins => fork92_outs_8,
      ins_valid => fork92_outs_8_valid,
      ins_ready => fork92_outs_8_ready,
      clk => clk,
      rst => rst,
      outs => buffer165_outs,
      outs_valid => buffer165_outs_valid,
      outs_ready => buffer165_outs_ready
    );

  sink19 : entity work.sink_dataless(arch)
    port map(
      ins_valid => cond_br129_falseOut_valid,
      ins_ready => cond_br129_falseOut_ready,
      clk => clk,
      rst => rst
    );

  cond_br130 : entity work.cond_br_dataless(arch)
    port map(
      condition => buffer166_outs,
      condition_valid => buffer166_outs_valid,
      condition_ready => buffer166_outs_ready,
      data_valid => fork76_outs_1_valid,
      data_ready => fork76_outs_1_ready,
      clk => clk,
      rst => rst,
      trueOut_valid => cond_br130_trueOut_valid,
      trueOut_ready => cond_br130_trueOut_ready,
      falseOut_valid => cond_br130_falseOut_valid,
      falseOut_ready => cond_br130_falseOut_ready
    );

  buffer166 : entity work.tfifo(arch) generic map(1, 1)
    port map(
      ins => fork92_outs_7,
      ins_valid => fork92_outs_7_valid,
      ins_ready => fork92_outs_7_ready,
      clk => clk,
      rst => rst,
      outs => buffer166_outs,
      outs_valid => buffer166_outs_valid,
      outs_ready => buffer166_outs_ready
    );

  sink20 : entity work.sink_dataless(arch)
    port map(
      ins_valid => cond_br130_falseOut_valid,
      ins_ready => cond_br130_falseOut_ready,
      clk => clk,
      rst => rst
    );

  cond_br131 : entity work.cond_br_dataless(arch)
    port map(
      condition => buffer167_outs,
      condition_valid => buffer167_outs_valid,
      condition_ready => buffer167_outs_ready,
      data_valid => fork78_outs_1_valid,
      data_ready => fork78_outs_1_ready,
      clk => clk,
      rst => rst,
      trueOut_valid => cond_br131_trueOut_valid,
      trueOut_ready => cond_br131_trueOut_ready,
      falseOut_valid => cond_br131_falseOut_valid,
      falseOut_ready => cond_br131_falseOut_ready
    );

  buffer167 : entity work.tfifo(arch) generic map(1, 1)
    port map(
      ins => fork92_outs_6,
      ins_valid => fork92_outs_6_valid,
      ins_ready => fork92_outs_6_ready,
      clk => clk,
      rst => rst,
      outs => buffer167_outs,
      outs_valid => buffer167_outs_valid,
      outs_ready => buffer167_outs_ready
    );

  sink21 : entity work.sink_dataless(arch)
    port map(
      ins_valid => cond_br131_falseOut_valid,
      ins_ready => cond_br131_falseOut_ready,
      clk => clk,
      rst => rst
    );

  cond_br132 : entity work.cond_br_dataless(arch)
    port map(
      condition => buffer168_outs,
      condition_valid => buffer168_outs_valid,
      condition_ready => buffer168_outs_ready,
      data_valid => buffer5_outs_valid,
      data_ready => buffer5_outs_ready,
      clk => clk,
      rst => rst,
      trueOut_valid => cond_br132_trueOut_valid,
      trueOut_ready => cond_br132_trueOut_ready,
      falseOut_valid => cond_br132_falseOut_valid,
      falseOut_ready => cond_br132_falseOut_ready
    );

  buffer168 : entity work.tfifo(arch) generic map(3, 1)
    port map(
      ins => fork92_outs_5,
      ins_valid => fork92_outs_5_valid,
      ins_ready => fork92_outs_5_ready,
      clk => clk,
      rst => rst,
      outs => buffer168_outs,
      outs_valid => buffer168_outs_valid,
      outs_ready => buffer168_outs_ready
    );

  cond_br133 : entity work.cond_br_dataless(arch)
    port map(
      condition => buffer169_outs,
      condition_valid => buffer169_outs_valid,
      condition_ready => buffer169_outs_ready,
      data_valid => fork77_outs_1_valid,
      data_ready => fork77_outs_1_ready,
      clk => clk,
      rst => rst,
      trueOut_valid => cond_br133_trueOut_valid,
      trueOut_ready => cond_br133_trueOut_ready,
      falseOut_valid => cond_br133_falseOut_valid,
      falseOut_ready => cond_br133_falseOut_ready
    );

  buffer169 : entity work.tfifo(arch) generic map(1, 1)
    port map(
      ins => fork92_outs_4,
      ins_valid => fork92_outs_4_valid,
      ins_ready => fork92_outs_4_ready,
      clk => clk,
      rst => rst,
      outs => buffer169_outs,
      outs_valid => buffer169_outs_valid,
      outs_ready => buffer169_outs_ready
    );

  sink22 : entity work.sink_dataless(arch)
    port map(
      ins_valid => cond_br133_falseOut_valid,
      ins_ready => cond_br133_falseOut_ready,
      clk => clk,
      rst => rst
    );

  init42 : entity work.tehb_init(arch) generic map(1, 0)
    port map(
      ins => fork92_outs_3,
      ins_valid => fork92_outs_3_valid,
      ins_ready => fork92_outs_3_ready,
      clk => clk,
      rst => rst,
      outs => init42_outs,
      outs_valid => init42_outs_valid,
      outs_ready => init42_outs_ready
    );

  fork74 : entity work.handshake_fork(arch) generic map(6, 1)
    port map(
      ins => init42_outs,
      ins_valid => init42_outs_valid,
      ins_ready => init42_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork74_outs_0,
      outs(1) => fork74_outs_1,
      outs(2) => fork74_outs_2,
      outs(3) => fork74_outs_3,
      outs(4) => fork74_outs_4,
      outs(5) => fork74_outs_5,
      outs_valid(0) => fork74_outs_0_valid,
      outs_valid(1) => fork74_outs_1_valid,
      outs_valid(2) => fork74_outs_2_valid,
      outs_valid(3) => fork74_outs_3_valid,
      outs_valid(4) => fork74_outs_4_valid,
      outs_valid(5) => fork74_outs_5_valid,
      outs_ready(0) => fork74_outs_0_ready,
      outs_ready(1) => fork74_outs_1_ready,
      outs_ready(2) => fork74_outs_2_ready,
      outs_ready(3) => fork74_outs_3_ready,
      outs_ready(4) => fork74_outs_4_ready,
      outs_ready(5) => fork74_outs_5_ready
    );

  mux60 : entity work.mux_dataless(arch) generic map(2, 1)
    port map(
      index => buffer171_outs,
      index_valid => buffer171_outs_valid,
      index_ready => buffer171_outs_ready,
      ins_valid(0) => buffer4_outs_valid,
      ins_valid(1) => cond_br129_trueOut_valid,
      ins_ready(0) => buffer4_outs_ready,
      ins_ready(1) => cond_br129_trueOut_ready,
      clk => clk,
      rst => rst,
      outs_valid => mux60_outs_valid,
      outs_ready => mux60_outs_ready
    );

  buffer171 : entity work.tfifo(arch) generic map(3, 1)
    port map(
      ins => fork74_outs_5,
      ins_valid => fork74_outs_5_valid,
      ins_ready => fork74_outs_5_ready,
      clk => clk,
      rst => rst,
      outs => buffer171_outs,
      outs_valid => buffer171_outs_valid,
      outs_ready => buffer171_outs_ready
    );

  buffer183 : entity work.oehb_dataless(arch)
    port map(
      ins_valid => mux60_outs_valid,
      ins_ready => mux60_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer183_outs_valid,
      outs_ready => buffer183_outs_ready
    );

  buffer184 : entity work.tehb_dataless(arch)
    port map(
      ins_valid => buffer183_outs_valid,
      ins_ready => buffer183_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer184_outs_valid,
      outs_ready => buffer184_outs_ready
    );

  fork75 : entity work.fork_dataless(arch) generic map(3)
    port map(
      ins_valid => buffer184_outs_valid,
      ins_ready => buffer184_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid(0) => fork75_outs_0_valid,
      outs_valid(1) => fork75_outs_1_valid,
      outs_valid(2) => fork75_outs_2_valid,
      outs_ready(0) => fork75_outs_0_ready,
      outs_ready(1) => fork75_outs_1_ready,
      outs_ready(2) => fork75_outs_2_ready
    );

  buffer180 : entity work.oehb_dataless(arch)
    port map(
      ins_valid => cond_br130_trueOut_valid,
      ins_ready => cond_br130_trueOut_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer180_outs_valid,
      outs_ready => buffer180_outs_ready
    );

  mux62 : entity work.mux_dataless(arch) generic map(2, 1)
    port map(
      index => buffer172_outs,
      index_valid => buffer172_outs_valid,
      index_ready => buffer172_outs_ready,
      ins_valid(0) => fork64_outs_1_valid,
      ins_valid(1) => buffer180_outs_valid,
      ins_ready(0) => fork64_outs_1_ready,
      ins_ready(1) => buffer180_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => mux62_outs_valid,
      outs_ready => mux62_outs_ready
    );

  buffer172 : entity work.tfifo(arch) generic map(1, 1)
    port map(
      ins => fork74_outs_4,
      ins_valid => fork74_outs_4_valid,
      ins_ready => fork74_outs_4_ready,
      clk => clk,
      rst => rst,
      outs => buffer172_outs,
      outs_valid => buffer172_outs_valid,
      outs_ready => buffer172_outs_ready
    );

  buffer186 : entity work.tehb_dataless(arch)
    port map(
      ins_valid => mux62_outs_valid,
      ins_ready => mux62_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer186_outs_valid,
      outs_ready => buffer186_outs_ready
    );

  fork76 : entity work.fork_dataless(arch) generic map(2)
    port map(
      ins_valid => buffer186_outs_valid,
      ins_ready => buffer186_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid(0) => fork76_outs_0_valid,
      outs_valid(1) => fork76_outs_1_valid,
      outs_ready(0) => fork76_outs_0_ready,
      outs_ready(1) => fork76_outs_1_ready
    );

  buffer182 : entity work.oehb_dataless(arch)
    port map(
      ins_valid => cond_br133_trueOut_valid,
      ins_ready => cond_br133_trueOut_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer182_outs_valid,
      outs_ready => buffer182_outs_ready
    );

  mux63 : entity work.mux_dataless(arch) generic map(2, 1)
    port map(
      index => buffer173_outs,
      index_valid => buffer173_outs_valid,
      index_ready => buffer173_outs_ready,
      ins_valid(0) => fork65_outs_1_valid,
      ins_valid(1) => buffer182_outs_valid,
      ins_ready(0) => fork65_outs_1_ready,
      ins_ready(1) => buffer182_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => mux63_outs_valid,
      outs_ready => mux63_outs_ready
    );

  buffer173 : entity work.tfifo(arch) generic map(1, 1)
    port map(
      ins => fork74_outs_3,
      ins_valid => fork74_outs_3_valid,
      ins_ready => fork74_outs_3_ready,
      clk => clk,
      rst => rst,
      outs => buffer173_outs,
      outs_valid => buffer173_outs_valid,
      outs_ready => buffer173_outs_ready
    );

  buffer188 : entity work.tehb_dataless(arch)
    port map(
      ins_valid => mux63_outs_valid,
      ins_ready => mux63_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer188_outs_valid,
      outs_ready => buffer188_outs_ready
    );

  fork77 : entity work.fork_dataless(arch) generic map(2)
    port map(
      ins_valid => buffer188_outs_valid,
      ins_ready => buffer188_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid(0) => fork77_outs_0_valid,
      outs_valid(1) => fork77_outs_1_valid,
      outs_ready(0) => fork77_outs_0_ready,
      outs_ready(1) => fork77_outs_1_ready
    );

  mux64 : entity work.mux_dataless(arch) generic map(2, 1)
    port map(
      index => buffer174_outs,
      index_valid => buffer174_outs_valid,
      index_ready => buffer174_outs_ready,
      ins_valid(0) => fork66_outs_1_valid,
      ins_valid(1) => cond_br131_trueOut_valid,
      ins_ready(0) => fork66_outs_1_ready,
      ins_ready(1) => cond_br131_trueOut_ready,
      clk => clk,
      rst => rst,
      outs_valid => mux64_outs_valid,
      outs_ready => mux64_outs_ready
    );

  buffer174 : entity work.tfifo(arch) generic map(1, 1)
    port map(
      ins => fork74_outs_2,
      ins_valid => fork74_outs_2_valid,
      ins_ready => fork74_outs_2_ready,
      clk => clk,
      rst => rst,
      outs => buffer174_outs,
      outs_valid => buffer174_outs_valid,
      outs_ready => buffer174_outs_ready
    );

  buffer191 : entity work.oehb_dataless(arch)
    port map(
      ins_valid => mux64_outs_valid,
      ins_ready => mux64_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer191_outs_valid,
      outs_ready => buffer191_outs_ready
    );

  buffer193 : entity work.tehb_dataless(arch)
    port map(
      ins_valid => buffer191_outs_valid,
      ins_ready => buffer191_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer193_outs_valid,
      outs_ready => buffer193_outs_ready
    );

  fork78 : entity work.fork_dataless(arch) generic map(2)
    port map(
      ins_valid => buffer193_outs_valid,
      ins_ready => buffer193_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid(0) => fork78_outs_0_valid,
      outs_valid(1) => fork78_outs_1_valid,
      outs_ready(0) => fork78_outs_0_ready,
      outs_ready(1) => fork78_outs_1_ready
    );

  mux65 : entity work.mux_dataless(arch) generic map(2, 1)
    port map(
      index => buffer175_outs,
      index_valid => buffer175_outs_valid,
      index_ready => buffer175_outs_ready,
      ins_valid(0) => fork67_outs_1_valid,
      ins_valid(1) => cond_br128_trueOut_valid,
      ins_ready(0) => fork67_outs_1_ready,
      ins_ready(1) => cond_br128_trueOut_ready,
      clk => clk,
      rst => rst,
      outs_valid => mux65_outs_valid,
      outs_ready => mux65_outs_ready
    );

  buffer175 : entity work.tfifo(arch) generic map(1, 1)
    port map(
      ins => fork74_outs_1,
      ins_valid => fork74_outs_1_valid,
      ins_ready => fork74_outs_1_ready,
      clk => clk,
      rst => rst,
      outs => buffer175_outs,
      outs_valid => buffer175_outs_valid,
      outs_ready => buffer175_outs_ready
    );

  buffer195 : entity work.tehb_dataless(arch)
    port map(
      ins_valid => mux65_outs_valid,
      ins_ready => mux65_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer195_outs_valid,
      outs_ready => buffer195_outs_ready
    );

  fork79 : entity work.fork_dataless(arch) generic map(2)
    port map(
      ins_valid => buffer195_outs_valid,
      ins_ready => buffer195_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid(0) => fork79_outs_0_valid,
      outs_valid(1) => fork79_outs_1_valid,
      outs_ready(0) => fork79_outs_0_ready,
      outs_ready(1) => fork79_outs_1_ready
    );

  buffer160 : entity work.tehb_dataless(arch)
    port map(
      ins_valid => mux58_outs_valid,
      ins_ready => mux58_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer160_outs_valid,
      outs_ready => buffer160_outs_ready
    );

  mux66 : entity work.mux_dataless(arch) generic map(2, 1)
    port map(
      index => buffer176_outs,
      index_valid => buffer176_outs_valid,
      index_ready => buffer176_outs_ready,
      ins_valid(0) => buffer160_outs_valid,
      ins_valid(1) => cond_br132_trueOut_valid,
      ins_ready(0) => buffer160_outs_ready,
      ins_ready(1) => cond_br132_trueOut_ready,
      clk => clk,
      rst => rst,
      outs_valid => mux66_outs_valid,
      outs_ready => mux66_outs_ready
    );

  buffer176 : entity work.tfifo(arch) generic map(3, 1)
    port map(
      ins => fork74_outs_0,
      ins_valid => fork74_outs_0_valid,
      ins_ready => fork74_outs_0_ready,
      clk => clk,
      rst => rst,
      outs => buffer176_outs,
      outs_valid => buffer176_outs_valid,
      outs_ready => buffer176_outs_ready
    );

  mux15 : entity work.mux(arch) generic map(2, 5, 1)
    port map(
      index => fork86_outs_2,
      index_valid => fork86_outs_2_valid,
      index_ready => fork86_outs_2_ready,
      ins(0) => extsi45_outs,
      ins(1) => cond_br29_trueOut,
      ins_valid(0) => extsi45_outs_valid,
      ins_valid(1) => cond_br29_trueOut_valid,
      ins_ready(0) => extsi45_outs_ready,
      ins_ready(1) => cond_br29_trueOut_ready,
      clk => clk,
      rst => rst,
      outs => mux15_outs,
      outs_valid => mux15_outs_valid,
      outs_ready => mux15_outs_ready
    );

  buffer215 : entity work.oehb(arch) generic map(5)
    port map(
      ins => mux15_outs,
      ins_valid => mux15_outs_valid,
      ins_ready => mux15_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer215_outs,
      outs_valid => buffer215_outs_valid,
      outs_ready => buffer215_outs_ready
    );

  buffer216 : entity work.tehb(arch) generic map(5)
    port map(
      ins => buffer215_outs,
      ins_valid => buffer215_outs_valid,
      ins_ready => buffer215_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer216_outs,
      outs_valid => buffer216_outs_valid,
      outs_ready => buffer216_outs_ready
    );

  fork80 : entity work.handshake_fork(arch) generic map(2, 5)
    port map(
      ins => buffer216_outs,
      ins_valid => buffer216_outs_valid,
      ins_ready => buffer216_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork80_outs_0,
      outs(1) => fork80_outs_1,
      outs_valid(0) => fork80_outs_0_valid,
      outs_valid(1) => fork80_outs_1_valid,
      outs_ready(0) => fork80_outs_0_ready,
      outs_ready(1) => fork80_outs_1_ready
    );

  extsi88 : entity work.extsi(arch) generic map(5, 6)
    port map(
      ins => fork80_outs_0,
      ins_valid => fork80_outs_0_valid,
      ins_ready => fork80_outs_0_ready,
      clk => clk,
      rst => rst,
      outs => extsi88_outs,
      outs_valid => extsi88_outs_valid,
      outs_ready => extsi88_outs_ready
    );

  extsi89 : entity work.extsi(arch) generic map(5, 32)
    port map(
      ins => fork80_outs_1,
      ins_valid => fork80_outs_1_valid,
      ins_ready => fork80_outs_1_ready,
      clk => clk,
      rst => rst,
      outs => extsi89_outs,
      outs_valid => extsi89_outs_valid,
      outs_ready => extsi89_outs_ready
    );

  fork81 : entity work.handshake_fork(arch) generic map(3, 32)
    port map(
      ins => extsi89_outs,
      ins_valid => extsi89_outs_valid,
      ins_ready => extsi89_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork81_outs_0,
      outs(1) => fork81_outs_1,
      outs(2) => fork81_outs_2,
      outs_valid(0) => fork81_outs_0_valid,
      outs_valid(1) => fork81_outs_1_valid,
      outs_valid(2) => fork81_outs_2_valid,
      outs_ready(0) => fork81_outs_0_ready,
      outs_ready(1) => fork81_outs_1_ready,
      outs_ready(2) => fork81_outs_2_ready
    );

  mux16 : entity work.mux(arch) generic map(2, 5, 1)
    port map(
      index => fork86_outs_0,
      index_valid => fork86_outs_0_valid,
      index_ready => fork86_outs_0_ready,
      ins(0) => fork69_outs_0,
      ins(1) => cond_br30_trueOut,
      ins_valid(0) => fork69_outs_0_valid,
      ins_valid(1) => cond_br30_trueOut_valid,
      ins_ready(0) => fork69_outs_0_ready,
      ins_ready(1) => cond_br30_trueOut_ready,
      clk => clk,
      rst => rst,
      outs => mux16_outs,
      outs_valid => mux16_outs_valid,
      outs_ready => mux16_outs_ready
    );

  buffer218 : entity work.oehb(arch) generic map(5)
    port map(
      ins => mux16_outs,
      ins_valid => mux16_outs_valid,
      ins_ready => mux16_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer218_outs,
      outs_valid => buffer218_outs_valid,
      outs_ready => buffer218_outs_ready
    );

  buffer220 : entity work.tehb(arch) generic map(5)
    port map(
      ins => buffer218_outs,
      ins_valid => buffer218_outs_valid,
      ins_ready => buffer218_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer220_outs,
      outs_valid => buffer220_outs_valid,
      outs_ready => buffer220_outs_ready
    );

  fork82 : entity work.handshake_fork(arch) generic map(2, 5)
    port map(
      ins => buffer220_outs,
      ins_valid => buffer220_outs_valid,
      ins_ready => buffer220_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork82_outs_0,
      outs(1) => fork82_outs_1,
      outs_valid(0) => fork82_outs_0_valid,
      outs_valid(1) => fork82_outs_1_valid,
      outs_ready(0) => fork82_outs_0_ready,
      outs_ready(1) => fork82_outs_1_ready
    );

  extsi90 : entity work.extsi(arch) generic map(5, 32)
    port map(
      ins => buffer181_outs,
      ins_valid => buffer181_outs_valid,
      ins_ready => buffer181_outs_ready,
      clk => clk,
      rst => rst,
      outs => extsi90_outs,
      outs_valid => extsi90_outs_valid,
      outs_ready => extsi90_outs_ready
    );

  buffer181 : entity work.tfifo(arch) generic map(1, 5)
    port map(
      ins => fork82_outs_1,
      ins_valid => fork82_outs_1_valid,
      ins_ready => fork82_outs_1_ready,
      clk => clk,
      rst => rst,
      outs => buffer181_outs,
      outs_valid => buffer181_outs_valid,
      outs_ready => buffer181_outs_ready
    );

  fork83 : entity work.handshake_fork(arch) generic map(6, 32)
    port map(
      ins => extsi90_outs,
      ins_valid => extsi90_outs_valid,
      ins_ready => extsi90_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork83_outs_0,
      outs(1) => fork83_outs_1,
      outs(2) => fork83_outs_2,
      outs(3) => fork83_outs_3,
      outs(4) => fork83_outs_4,
      outs(5) => fork83_outs_5,
      outs_valid(0) => fork83_outs_0_valid,
      outs_valid(1) => fork83_outs_1_valid,
      outs_valid(2) => fork83_outs_2_valid,
      outs_valid(3) => fork83_outs_3_valid,
      outs_valid(4) => fork83_outs_4_valid,
      outs_valid(5) => fork83_outs_5_valid,
      outs_ready(0) => fork83_outs_0_ready,
      outs_ready(1) => fork83_outs_1_ready,
      outs_ready(2) => fork83_outs_2_ready,
      outs_ready(3) => fork83_outs_3_ready,
      outs_ready(4) => fork83_outs_4_ready,
      outs_ready(5) => fork83_outs_5_ready
    );

  mux17 : entity work.mux(arch) generic map(2, 5, 1)
    port map(
      index => fork86_outs_1,
      index_valid => fork86_outs_1_valid,
      index_ready => fork86_outs_1_ready,
      ins(0) => fork68_outs_1,
      ins(1) => cond_br31_trueOut,
      ins_valid(0) => fork68_outs_1_valid,
      ins_valid(1) => cond_br31_trueOut_valid,
      ins_ready(0) => fork68_outs_1_ready,
      ins_ready(1) => cond_br31_trueOut_ready,
      clk => clk,
      rst => rst,
      outs => mux17_outs,
      outs_valid => mux17_outs_valid,
      outs_ready => mux17_outs_ready
    );

  buffer221 : entity work.oehb(arch) generic map(5)
    port map(
      ins => mux17_outs,
      ins_valid => mux17_outs_valid,
      ins_ready => mux17_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer221_outs,
      outs_valid => buffer221_outs_valid,
      outs_ready => buffer221_outs_ready
    );

  buffer222 : entity work.tehb(arch) generic map(5)
    port map(
      ins => buffer221_outs,
      ins_valid => buffer221_outs_valid,
      ins_ready => buffer221_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer222_outs,
      outs_valid => buffer222_outs_valid,
      outs_ready => buffer222_outs_ready
    );

  fork84 : entity work.handshake_fork(arch) generic map(2, 5)
    port map(
      ins => buffer222_outs,
      ins_valid => buffer222_outs_valid,
      ins_ready => buffer222_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork84_outs_0,
      outs(1) => fork84_outs_1,
      outs_valid(0) => fork84_outs_0_valid,
      outs_valid(1) => fork84_outs_1_valid,
      outs_ready(0) => fork84_outs_0_ready,
      outs_ready(1) => fork84_outs_1_ready
    );

  extsi91 : entity work.extsi(arch) generic map(5, 32)
    port map(
      ins => fork84_outs_1,
      ins_valid => fork84_outs_1_valid,
      ins_ready => fork84_outs_1_ready,
      clk => clk,
      rst => rst,
      outs => extsi91_outs,
      outs_valid => extsi91_outs_valid,
      outs_ready => extsi91_outs_ready
    );

  fork85 : entity work.handshake_fork(arch) generic map(3, 32)
    port map(
      ins => extsi91_outs,
      ins_valid => extsi91_outs_valid,
      ins_ready => extsi91_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork85_outs_0,
      outs(1) => fork85_outs_1,
      outs(2) => fork85_outs_2,
      outs_valid(0) => fork85_outs_0_valid,
      outs_valid(1) => fork85_outs_1_valid,
      outs_valid(2) => fork85_outs_2_valid,
      outs_ready(0) => fork85_outs_0_ready,
      outs_ready(1) => fork85_outs_1_ready,
      outs_ready(2) => fork85_outs_2_ready
    );

  control_merge12 : entity work.control_merge_dataless(arch) generic map(2, 1)
    port map(
      ins_valid(0) => fork72_outs_2_valid,
      ins_valid(1) => cond_br32_trueOut_valid,
      ins_ready(0) => fork72_outs_2_ready,
      ins_ready(1) => cond_br32_trueOut_ready,
      clk => clk,
      rst => rst,
      outs_valid => control_merge12_outs_valid,
      outs_ready => control_merge12_outs_ready,
      index => control_merge12_index,
      index_valid => control_merge12_index_valid,
      index_ready => control_merge12_index_ready
    );

  fork86 : entity work.handshake_fork(arch) generic map(3, 1)
    port map(
      ins => control_merge12_index,
      ins_valid => control_merge12_index_valid,
      ins_ready => control_merge12_index_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork86_outs_0,
      outs(1) => fork86_outs_1,
      outs(2) => fork86_outs_2,
      outs_valid(0) => fork86_outs_0_valid,
      outs_valid(1) => fork86_outs_1_valid,
      outs_valid(2) => fork86_outs_2_valid,
      outs_ready(0) => fork86_outs_0_ready,
      outs_ready(1) => fork86_outs_1_ready,
      outs_ready(2) => fork86_outs_2_ready
    );

  buffer224 : entity work.oehb_dataless(arch)
    port map(
      ins_valid => control_merge12_outs_valid,
      ins_ready => control_merge12_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer224_outs_valid,
      outs_ready => buffer224_outs_ready
    );

  fork87 : entity work.fork_dataless(arch) generic map(2)
    port map(
      ins_valid => buffer224_outs_valid,
      ins_ready => buffer224_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid(0) => fork87_outs_0_valid,
      outs_valid(1) => fork87_outs_1_valid,
      outs_ready(0) => fork87_outs_0_ready,
      outs_ready(1) => fork87_outs_1_ready
    );

  constant79 : entity work.handshake_constant_1(arch) generic map(2)
    port map(
      ctrl_valid => fork87_outs_0_valid,
      ctrl_ready => fork87_outs_0_ready,
      clk => clk,
      rst => rst,
      outs => constant79_outs,
      outs_valid => constant79_outs_valid,
      outs_ready => constant79_outs_ready
    );

  extsi37 : entity work.extsi(arch) generic map(2, 32)
    port map(
      ins => constant79_outs,
      ins_valid => constant79_outs_valid,
      ins_ready => constant79_outs_ready,
      clk => clk,
      rst => rst,
      outs => extsi37_outs,
      outs_valid => extsi37_outs_valid,
      outs_ready => extsi37_outs_ready
    );

  source20 : entity work.source(arch)
    port map(
      clk => clk,
      rst => rst,
      outs_valid => source20_outs_valid,
      outs_ready => source20_outs_ready
    );

  constant80 : entity work.handshake_constant_3(arch) generic map(5)
    port map(
      ctrl_valid => source20_outs_valid,
      ctrl_ready => source20_outs_ready,
      clk => clk,
      rst => rst,
      outs => constant80_outs,
      outs_valid => constant80_outs_valid,
      outs_ready => constant80_outs_ready
    );

  extsi92 : entity work.extsi(arch) generic map(5, 6)
    port map(
      ins => constant80_outs,
      ins_valid => constant80_outs_valid,
      ins_ready => constant80_outs_ready,
      clk => clk,
      rst => rst,
      outs => extsi92_outs,
      outs_valid => extsi92_outs_valid,
      outs_ready => extsi92_outs_ready
    );

  source21 : entity work.source(arch)
    port map(
      clk => clk,
      rst => rst,
      outs_valid => source21_outs_valid,
      outs_ready => source21_outs_ready
    );

  constant81 : entity work.handshake_constant_1(arch) generic map(2)
    port map(
      ctrl_valid => source21_outs_valid,
      ctrl_ready => source21_outs_ready,
      clk => clk,
      rst => rst,
      outs => constant81_outs,
      outs_valid => constant81_outs_valid,
      outs_ready => constant81_outs_ready
    );

  fork88 : entity work.handshake_fork(arch) generic map(2, 2)
    port map(
      ins => constant81_outs,
      ins_valid => constant81_outs_valid,
      ins_ready => constant81_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork88_outs_0,
      outs(1) => fork88_outs_1,
      outs_valid(0) => fork88_outs_0_valid,
      outs_valid(1) => fork88_outs_1_valid,
      outs_ready(0) => fork88_outs_0_ready,
      outs_ready(1) => fork88_outs_1_ready
    );

  extsi93 : entity work.extsi(arch) generic map(2, 6)
    port map(
      ins => fork88_outs_0,
      ins_valid => fork88_outs_0_valid,
      ins_ready => fork88_outs_0_ready,
      clk => clk,
      rst => rst,
      outs => extsi93_outs,
      outs_valid => extsi93_outs_valid,
      outs_ready => extsi93_outs_ready
    );

  extsi39 : entity work.extsi(arch) generic map(2, 32)
    port map(
      ins => buffer185_outs,
      ins_valid => buffer185_outs_valid,
      ins_ready => buffer185_outs_ready,
      clk => clk,
      rst => rst,
      outs => extsi39_outs,
      outs_valid => extsi39_outs_valid,
      outs_ready => extsi39_outs_ready
    );

  buffer185 : entity work.tfifo(arch) generic map(1, 2)
    port map(
      ins => fork88_outs_1,
      ins_valid => fork88_outs_1_valid,
      ins_ready => fork88_outs_1_ready,
      clk => clk,
      rst => rst,
      outs => buffer185_outs,
      outs_valid => buffer185_outs_valid,
      outs_ready => buffer185_outs_ready
    );

  fork89 : entity work.handshake_fork(arch) generic map(4, 32)
    port map(
      ins => extsi39_outs,
      ins_valid => extsi39_outs_valid,
      ins_ready => extsi39_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork89_outs_0,
      outs(1) => fork89_outs_1,
      outs(2) => fork89_outs_2,
      outs(3) => fork89_outs_3,
      outs_valid(0) => fork89_outs_0_valid,
      outs_valid(1) => fork89_outs_1_valid,
      outs_valid(2) => fork89_outs_2_valid,
      outs_valid(3) => fork89_outs_3_valid,
      outs_ready(0) => fork89_outs_0_ready,
      outs_ready(1) => fork89_outs_1_ready,
      outs_ready(2) => fork89_outs_2_ready,
      outs_ready(3) => fork89_outs_3_ready
    );

  source22 : entity work.source(arch)
    port map(
      clk => clk,
      rst => rst,
      outs_valid => source22_outs_valid,
      outs_ready => source22_outs_ready
    );

  constant82 : entity work.handshake_constant_2(arch) generic map(3)
    port map(
      ctrl_valid => source22_outs_valid,
      ctrl_ready => source22_outs_ready,
      clk => clk,
      rst => rst,
      outs => constant82_outs,
      outs_valid => constant82_outs_valid,
      outs_ready => constant82_outs_ready
    );

  extsi40 : entity work.extsi(arch) generic map(3, 32)
    port map(
      ins => constant82_outs,
      ins_valid => constant82_outs_valid,
      ins_ready => constant82_outs_ready,
      clk => clk,
      rst => rst,
      outs => extsi40_outs,
      outs_valid => extsi40_outs_valid,
      outs_ready => extsi40_outs_ready
    );

  fork90 : entity work.handshake_fork(arch) generic map(4, 32)
    port map(
      ins => extsi40_outs,
      ins_valid => extsi40_outs_valid,
      ins_ready => extsi40_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork90_outs_0,
      outs(1) => fork90_outs_1,
      outs(2) => fork90_outs_2,
      outs(3) => fork90_outs_3,
      outs_valid(0) => fork90_outs_0_valid,
      outs_valid(1) => fork90_outs_1_valid,
      outs_valid(2) => fork90_outs_2_valid,
      outs_valid(3) => fork90_outs_3_valid,
      outs_ready(0) => fork90_outs_0_ready,
      outs_ready(1) => fork90_outs_1_ready,
      outs_ready(2) => fork90_outs_2_ready,
      outs_ready(3) => fork90_outs_3_ready
    );

  shli22 : entity work.shli(arch) generic map(32)
    port map(
      lhs => buffer187_outs,
      lhs_valid => buffer187_outs_valid,
      lhs_ready => buffer187_outs_ready,
      rhs => fork89_outs_0,
      rhs_valid => fork89_outs_0_valid,
      rhs_ready => fork89_outs_0_ready,
      clk => clk,
      rst => rst,
      result => shli22_result,
      result_valid => shli22_result_valid,
      result_ready => shli22_result_ready
    );

  buffer187 : entity work.tfifo(arch) generic map(1, 32)
    port map(
      ins => fork83_outs_0,
      ins_valid => fork83_outs_0_valid,
      ins_ready => fork83_outs_0_ready,
      clk => clk,
      rst => rst,
      outs => buffer187_outs,
      outs_valid => buffer187_outs_valid,
      outs_ready => buffer187_outs_ready
    );

  shli23 : entity work.shli(arch) generic map(32)
    port map(
      lhs => buffer189_outs,
      lhs_valid => buffer189_outs_valid,
      lhs_ready => buffer189_outs_ready,
      rhs => fork90_outs_0,
      rhs_valid => fork90_outs_0_valid,
      rhs_ready => fork90_outs_0_ready,
      clk => clk,
      rst => rst,
      result => shli23_result,
      result_valid => shli23_result_valid,
      result_ready => shli23_result_ready
    );

  buffer189 : entity work.tfifo(arch) generic map(1, 32)
    port map(
      ins => fork83_outs_1,
      ins_valid => fork83_outs_1_valid,
      ins_ready => fork83_outs_1_ready,
      clk => clk,
      rst => rst,
      outs => buffer189_outs,
      outs_valid => buffer189_outs_valid,
      outs_ready => buffer189_outs_ready
    );

  buffer226 : entity work.oehb(arch) generic map(32)
    port map(
      ins => shli22_result,
      ins_valid => shli22_result_valid,
      ins_ready => shli22_result_ready,
      clk => clk,
      rst => rst,
      outs => buffer226_outs,
      outs_valid => buffer226_outs_valid,
      outs_ready => buffer226_outs_ready
    );

  buffer227 : entity work.oehb(arch) generic map(32)
    port map(
      ins => shli23_result,
      ins_valid => shli23_result_valid,
      ins_ready => shli23_result_ready,
      clk => clk,
      rst => rst,
      outs => buffer227_outs,
      outs_valid => buffer227_outs_valid,
      outs_ready => buffer227_outs_ready
    );

  addi38 : entity work.addi(arch) generic map(32)
    port map(
      lhs => buffer226_outs,
      lhs_valid => buffer226_outs_valid,
      lhs_ready => buffer226_outs_ready,
      rhs => buffer227_outs,
      rhs_valid => buffer227_outs_valid,
      rhs_ready => buffer227_outs_ready,
      clk => clk,
      rst => rst,
      result => addi38_result,
      result_valid => addi38_result_valid,
      result_ready => addi38_result_ready
    );

  buffer228 : entity work.oehb(arch) generic map(32)
    port map(
      ins => addi38_result,
      ins_valid => addi38_result_valid,
      ins_ready => addi38_result_ready,
      clk => clk,
      rst => rst,
      outs => buffer228_outs,
      outs_valid => buffer228_outs_valid,
      outs_ready => buffer228_outs_ready
    );

  addi14 : entity work.addi(arch) generic map(32)
    port map(
      lhs => buffer190_outs,
      lhs_valid => buffer190_outs_valid,
      lhs_ready => buffer190_outs_ready,
      rhs => buffer228_outs,
      rhs_valid => buffer228_outs_valid,
      rhs_ready => buffer228_outs_ready,
      clk => clk,
      rst => rst,
      result => addi14_result,
      result_valid => addi14_result_valid,
      result_ready => addi14_result_ready
    );

  buffer190 : entity work.tfifo(arch) generic map(1, 32)
    port map(
      ins => fork81_outs_0,
      ins_valid => fork81_outs_0_valid,
      ins_ready => fork81_outs_0_ready,
      clk => clk,
      rst => rst,
      outs => buffer190_outs,
      outs_valid => buffer190_outs_valid,
      outs_ready => buffer190_outs_ready
    );

  gate4 : entity work.gate(arch) generic map(3, 32)
    port map(
      ins(0) => addi14_result,
      ins_valid(0) => addi14_result_valid,
      ins_valid(1) => fork79_outs_0_valid,
      ins_valid(2) => fork78_outs_0_valid,
      ins_ready(0) => addi14_result_ready,
      ins_ready(1) => fork79_outs_0_ready,
      ins_ready(2) => fork78_outs_0_ready,
      clk => clk,
      rst => rst,
      outs => gate4_outs,
      outs_valid => gate4_outs_valid,
      outs_ready => gate4_outs_ready
    );

  trunci24 : entity work.trunci(arch) generic map(32, 7)
    port map(
      ins => gate4_outs,
      ins_valid => gate4_outs_valid,
      ins_ready => gate4_outs_ready,
      clk => clk,
      rst => rst,
      outs => trunci24_outs,
      outs_valid => trunci24_outs_valid,
      outs_ready => trunci24_outs_ready
    );

  load6 : entity work.load(arch) generic map(32, 7)
    port map(
      addrIn => trunci24_outs,
      addrIn_valid => trunci24_outs_valid,
      addrIn_ready => trunci24_outs_ready,
      dataFromMem => mem_controller6_ldData_1,
      dataFromMem_valid => mem_controller6_ldData_1_valid,
      dataFromMem_ready => mem_controller6_ldData_1_ready,
      clk => clk,
      rst => rst,
      addrOut => load6_addrOut,
      addrOut_valid => load6_addrOut_valid,
      addrOut_ready => load6_addrOut_ready,
      dataOut => load6_dataOut,
      dataOut_valid => load6_dataOut_valid,
      dataOut_ready => load6_dataOut_ready
    );

  shli24 : entity work.shli(arch) generic map(32)
    port map(
      lhs => buffer192_outs,
      lhs_valid => buffer192_outs_valid,
      lhs_ready => buffer192_outs_ready,
      rhs => fork89_outs_1,
      rhs_valid => fork89_outs_1_valid,
      rhs_ready => fork89_outs_1_ready,
      clk => clk,
      rst => rst,
      result => shli24_result,
      result_valid => shli24_result_valid,
      result_ready => shli24_result_ready
    );

  buffer192 : entity work.tfifo(arch) generic map(1, 32)
    port map(
      ins => fork81_outs_1,
      ins_valid => fork81_outs_1_valid,
      ins_ready => fork81_outs_1_ready,
      clk => clk,
      rst => rst,
      outs => buffer192_outs,
      outs_valid => buffer192_outs_valid,
      outs_ready => buffer192_outs_ready
    );

  shli25 : entity work.shli(arch) generic map(32)
    port map(
      lhs => buffer194_outs,
      lhs_valid => buffer194_outs_valid,
      lhs_ready => buffer194_outs_ready,
      rhs => fork90_outs_1,
      rhs_valid => fork90_outs_1_valid,
      rhs_ready => fork90_outs_1_ready,
      clk => clk,
      rst => rst,
      result => shli25_result,
      result_valid => shli25_result_valid,
      result_ready => shli25_result_ready
    );

  buffer194 : entity work.tfifo(arch) generic map(1, 32)
    port map(
      ins => fork81_outs_2,
      ins_valid => fork81_outs_2_valid,
      ins_ready => fork81_outs_2_ready,
      clk => clk,
      rst => rst,
      outs => buffer194_outs,
      outs_valid => buffer194_outs_valid,
      outs_ready => buffer194_outs_ready
    );

  buffer229 : entity work.oehb(arch) generic map(32)
    port map(
      ins => shli24_result,
      ins_valid => shli24_result_valid,
      ins_ready => shli24_result_ready,
      clk => clk,
      rst => rst,
      outs => buffer229_outs,
      outs_valid => buffer229_outs_valid,
      outs_ready => buffer229_outs_ready
    );

  buffer230 : entity work.oehb(arch) generic map(32)
    port map(
      ins => shli25_result,
      ins_valid => shli25_result_valid,
      ins_ready => shli25_result_ready,
      clk => clk,
      rst => rst,
      outs => buffer230_outs,
      outs_valid => buffer230_outs_valid,
      outs_ready => buffer230_outs_ready
    );

  addi39 : entity work.addi(arch) generic map(32)
    port map(
      lhs => buffer229_outs,
      lhs_valid => buffer229_outs_valid,
      lhs_ready => buffer229_outs_ready,
      rhs => buffer230_outs,
      rhs_valid => buffer230_outs_valid,
      rhs_ready => buffer230_outs_ready,
      clk => clk,
      rst => rst,
      result => addi39_result,
      result_valid => addi39_result_valid,
      result_ready => addi39_result_ready
    );

  buffer231 : entity work.oehb(arch) generic map(32)
    port map(
      ins => addi39_result,
      ins_valid => addi39_result_valid,
      ins_ready => addi39_result_ready,
      clk => clk,
      rst => rst,
      outs => buffer231_outs,
      outs_valid => buffer231_outs_valid,
      outs_ready => buffer231_outs_ready
    );

  addi15 : entity work.addi(arch) generic map(32)
    port map(
      lhs => fork85_outs_0,
      lhs_valid => fork85_outs_0_valid,
      lhs_ready => fork85_outs_0_ready,
      rhs => buffer231_outs,
      rhs_valid => buffer231_outs_valid,
      rhs_ready => buffer231_outs_ready,
      clk => clk,
      rst => rst,
      result => addi15_result,
      result_valid => addi15_result_valid,
      result_ready => addi15_result_ready
    );

  gate5 : entity work.gate(arch) generic map(3, 32)
    port map(
      ins(0) => addi15_result,
      ins_valid(0) => addi15_result_valid,
      ins_valid(1) => fork77_outs_0_valid,
      ins_valid(2) => fork76_outs_0_valid,
      ins_ready(0) => addi15_result_ready,
      ins_ready(1) => fork77_outs_0_ready,
      ins_ready(2) => fork76_outs_0_ready,
      clk => clk,
      rst => rst,
      outs => gate5_outs,
      outs_valid => gate5_outs_valid,
      outs_ready => gate5_outs_ready
    );

  trunci25 : entity work.trunci(arch) generic map(32, 7)
    port map(
      ins => gate5_outs,
      ins_valid => gate5_outs_valid,
      ins_ready => gate5_outs_ready,
      clk => clk,
      rst => rst,
      outs => trunci25_outs,
      outs_valid => trunci25_outs_valid,
      outs_ready => trunci25_outs_ready
    );

  load7 : entity work.load(arch) generic map(32, 7)
    port map(
      addrIn => trunci25_outs,
      addrIn_valid => trunci25_outs_valid,
      addrIn_ready => trunci25_outs_ready,
      dataFromMem => mem_controller5_ldData_1,
      dataFromMem_valid => mem_controller5_ldData_1_valid,
      dataFromMem_ready => mem_controller5_ldData_1_ready,
      clk => clk,
      rst => rst,
      addrOut => load7_addrOut,
      addrOut_valid => load7_addrOut_valid,
      addrOut_ready => load7_addrOut_ready,
      dataOut => load7_dataOut,
      dataOut_valid => load7_dataOut_valid,
      dataOut_ready => load7_dataOut_ready
    );

  muli2 : entity work.muli(arch) generic map(32)
    port map(
      lhs => load6_dataOut,
      lhs_valid => load6_dataOut_valid,
      lhs_ready => load6_dataOut_ready,
      rhs => load7_dataOut,
      rhs_valid => load7_dataOut_valid,
      rhs_ready => load7_dataOut_ready,
      clk => clk,
      rst => rst,
      result => muli2_result,
      result_valid => muli2_result_valid,
      result_ready => muli2_result_ready
    );

  shli26 : entity work.shli(arch) generic map(32)
    port map(
      lhs => buffer197_outs,
      lhs_valid => buffer197_outs_valid,
      lhs_ready => buffer197_outs_ready,
      rhs => buffer196_outs,
      rhs_valid => buffer196_outs_valid,
      rhs_ready => buffer196_outs_ready,
      clk => clk,
      rst => rst,
      result => shli26_result,
      result_valid => shli26_result_valid,
      result_ready => shli26_result_ready
    );

  buffer196 : entity work.tfifo(arch) generic map(3, 32)
    port map(
      ins => fork89_outs_2,
      ins_valid => fork89_outs_2_valid,
      ins_ready => fork89_outs_2_ready,
      clk => clk,
      rst => rst,
      outs => buffer196_outs,
      outs_valid => buffer196_outs_valid,
      outs_ready => buffer196_outs_ready
    );

  buffer197 : entity work.tfifo(arch) generic map(2, 32)
    port map(
      ins => fork83_outs_2,
      ins_valid => fork83_outs_2_valid,
      ins_ready => fork83_outs_2_ready,
      clk => clk,
      rst => rst,
      outs => buffer197_outs,
      outs_valid => buffer197_outs_valid,
      outs_ready => buffer197_outs_ready
    );

  shli27 : entity work.shli(arch) generic map(32)
    port map(
      lhs => buffer199_outs,
      lhs_valid => buffer199_outs_valid,
      lhs_ready => buffer199_outs_ready,
      rhs => buffer198_outs,
      rhs_valid => buffer198_outs_valid,
      rhs_ready => buffer198_outs_ready,
      clk => clk,
      rst => rst,
      result => shli27_result,
      result_valid => shli27_result_valid,
      result_ready => shli27_result_ready
    );

  buffer198 : entity work.tfifo(arch) generic map(3, 32)
    port map(
      ins => fork90_outs_2,
      ins_valid => fork90_outs_2_valid,
      ins_ready => fork90_outs_2_ready,
      clk => clk,
      rst => rst,
      outs => buffer198_outs,
      outs_valid => buffer198_outs_valid,
      outs_ready => buffer198_outs_ready
    );

  buffer199 : entity work.tfifo(arch) generic map(2, 32)
    port map(
      ins => fork83_outs_3,
      ins_valid => fork83_outs_3_valid,
      ins_ready => fork83_outs_3_ready,
      clk => clk,
      rst => rst,
      outs => buffer199_outs,
      outs_valid => buffer199_outs_valid,
      outs_ready => buffer199_outs_ready
    );

  buffer233 : entity work.oehb(arch) generic map(32)
    port map(
      ins => shli26_result,
      ins_valid => shli26_result_valid,
      ins_ready => shli26_result_ready,
      clk => clk,
      rst => rst,
      outs => buffer233_outs,
      outs_valid => buffer233_outs_valid,
      outs_ready => buffer233_outs_ready
    );

  buffer234 : entity work.oehb(arch) generic map(32)
    port map(
      ins => shli27_result,
      ins_valid => shli27_result_valid,
      ins_ready => shli27_result_ready,
      clk => clk,
      rst => rst,
      outs => buffer234_outs,
      outs_valid => buffer234_outs_valid,
      outs_ready => buffer234_outs_ready
    );

  addi40 : entity work.addi(arch) generic map(32)
    port map(
      lhs => buffer233_outs,
      lhs_valid => buffer233_outs_valid,
      lhs_ready => buffer233_outs_ready,
      rhs => buffer234_outs,
      rhs_valid => buffer234_outs_valid,
      rhs_ready => buffer234_outs_ready,
      clk => clk,
      rst => rst,
      result => addi40_result,
      result_valid => addi40_result_valid,
      result_ready => addi40_result_ready
    );

  buffer235 : entity work.oehb(arch) generic map(32)
    port map(
      ins => addi40_result,
      ins_valid => addi40_result_valid,
      ins_ready => addi40_result_ready,
      clk => clk,
      rst => rst,
      outs => buffer235_outs,
      outs_valid => buffer235_outs_valid,
      outs_ready => buffer235_outs_ready
    );

  addi16 : entity work.addi(arch) generic map(32)
    port map(
      lhs => buffer200_outs,
      lhs_valid => buffer200_outs_valid,
      lhs_ready => buffer200_outs_ready,
      rhs => buffer235_outs,
      rhs_valid => buffer235_outs_valid,
      rhs_ready => buffer235_outs_ready,
      clk => clk,
      rst => rst,
      result => addi16_result,
      result_valid => addi16_result_valid,
      result_ready => addi16_result_ready
    );

  buffer200 : entity work.tfifo(arch) generic map(2, 32)
    port map(
      ins => fork85_outs_1,
      ins_valid => fork85_outs_1_valid,
      ins_ready => fork85_outs_1_ready,
      clk => clk,
      rst => rst,
      outs => buffer200_outs,
      outs_valid => buffer200_outs_valid,
      outs_ready => buffer200_outs_ready
    );

  buffer211 : entity work.tehb_dataless(arch)
    port map(
      ins_valid => mux66_outs_valid,
      ins_ready => mux66_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer211_outs_valid,
      outs_ready => buffer211_outs_ready
    );

  gate6 : entity work.gate(arch) generic map(3, 32)
    port map(
      ins(0) => addi16_result,
      ins_valid(0) => addi16_result_valid,
      ins_valid(1) => fork75_outs_1_valid,
      ins_valid(2) => buffer211_outs_valid,
      ins_ready(0) => addi16_result_ready,
      ins_ready(1) => fork75_outs_1_ready,
      ins_ready(2) => buffer211_outs_ready,
      clk => clk,
      rst => rst,
      outs => gate6_outs,
      outs_valid => gate6_outs_valid,
      outs_ready => gate6_outs_ready
    );

  trunci26 : entity work.trunci(arch) generic map(32, 7)
    port map(
      ins => gate6_outs,
      ins_valid => gate6_outs_valid,
      ins_ready => gate6_outs_ready,
      clk => clk,
      rst => rst,
      outs => trunci26_outs,
      outs_valid => trunci26_outs_valid,
      outs_ready => trunci26_outs_ready
    );

  load8 : entity work.load(arch) generic map(32, 7)
    port map(
      addrIn => trunci26_outs,
      addrIn_valid => trunci26_outs_valid,
      addrIn_ready => trunci26_outs_ready,
      dataFromMem => mem_controller4_ldData_0,
      dataFromMem_valid => mem_controller4_ldData_0_valid,
      dataFromMem_ready => mem_controller4_ldData_0_ready,
      clk => clk,
      rst => rst,
      addrOut => load8_addrOut,
      addrOut_valid => load8_addrOut_valid,
      addrOut_ready => load8_addrOut_ready,
      dataOut => load8_dataOut,
      dataOut_valid => load8_dataOut_valid,
      dataOut_ready => load8_dataOut_ready
    );

  addi2 : entity work.addi(arch) generic map(32)
    port map(
      lhs => load8_dataOut,
      lhs_valid => load8_dataOut_valid,
      lhs_ready => load8_dataOut_ready,
      rhs => muli2_result,
      rhs_valid => muli2_result_valid,
      rhs_ready => muli2_result_ready,
      clk => clk,
      rst => rst,
      result => addi2_result,
      result_valid => addi2_result_valid,
      result_ready => addi2_result_ready
    );

  shli28 : entity work.shli(arch) generic map(32)
    port map(
      lhs => buffer202_outs,
      lhs_valid => buffer202_outs_valid,
      lhs_ready => buffer202_outs_ready,
      rhs => buffer201_outs,
      rhs_valid => buffer201_outs_valid,
      rhs_ready => buffer201_outs_ready,
      clk => clk,
      rst => rst,
      result => shli28_result,
      result_valid => shli28_result_valid,
      result_ready => shli28_result_ready
    );

  buffer201 : entity work.tfifo(arch) generic map(2, 32)
    port map(
      ins => fork89_outs_3,
      ins_valid => fork89_outs_3_valid,
      ins_ready => fork89_outs_3_ready,
      clk => clk,
      rst => rst,
      outs => buffer201_outs,
      outs_valid => buffer201_outs_valid,
      outs_ready => buffer201_outs_ready
    );

  buffer202 : entity work.tfifo(arch) generic map(2, 32)
    port map(
      ins => fork83_outs_4,
      ins_valid => fork83_outs_4_valid,
      ins_ready => fork83_outs_4_ready,
      clk => clk,
      rst => rst,
      outs => buffer202_outs,
      outs_valid => buffer202_outs_valid,
      outs_ready => buffer202_outs_ready
    );

  shli29 : entity work.shli(arch) generic map(32)
    port map(
      lhs => buffer204_outs,
      lhs_valid => buffer204_outs_valid,
      lhs_ready => buffer204_outs_ready,
      rhs => buffer203_outs,
      rhs_valid => buffer203_outs_valid,
      rhs_ready => buffer203_outs_ready,
      clk => clk,
      rst => rst,
      result => shli29_result,
      result_valid => shli29_result_valid,
      result_ready => shli29_result_ready
    );

  buffer203 : entity work.tfifo(arch) generic map(2, 32)
    port map(
      ins => fork90_outs_3,
      ins_valid => fork90_outs_3_valid,
      ins_ready => fork90_outs_3_ready,
      clk => clk,
      rst => rst,
      outs => buffer203_outs,
      outs_valid => buffer203_outs_valid,
      outs_ready => buffer203_outs_ready
    );

  buffer204 : entity work.tfifo(arch) generic map(2, 32)
    port map(
      ins => fork83_outs_5,
      ins_valid => fork83_outs_5_valid,
      ins_ready => fork83_outs_5_ready,
      clk => clk,
      rst => rst,
      outs => buffer204_outs,
      outs_valid => buffer204_outs_valid,
      outs_ready => buffer204_outs_ready
    );

  buffer236 : entity work.oehb(arch) generic map(32)
    port map(
      ins => shli28_result,
      ins_valid => shli28_result_valid,
      ins_ready => shli28_result_ready,
      clk => clk,
      rst => rst,
      outs => buffer236_outs,
      outs_valid => buffer236_outs_valid,
      outs_ready => buffer236_outs_ready
    );

  buffer237 : entity work.oehb(arch) generic map(32)
    port map(
      ins => shli29_result,
      ins_valid => shli29_result_valid,
      ins_ready => shli29_result_ready,
      clk => clk,
      rst => rst,
      outs => buffer237_outs,
      outs_valid => buffer237_outs_valid,
      outs_ready => buffer237_outs_ready
    );

  addi41 : entity work.addi(arch) generic map(32)
    port map(
      lhs => buffer236_outs,
      lhs_valid => buffer236_outs_valid,
      lhs_ready => buffer236_outs_ready,
      rhs => buffer237_outs,
      rhs_valid => buffer237_outs_valid,
      rhs_ready => buffer237_outs_ready,
      clk => clk,
      rst => rst,
      result => addi41_result,
      result_valid => addi41_result_valid,
      result_ready => addi41_result_ready
    );

  buffer238 : entity work.oehb(arch) generic map(32)
    port map(
      ins => addi41_result,
      ins_valid => addi41_result_valid,
      ins_ready => addi41_result_ready,
      clk => clk,
      rst => rst,
      outs => buffer238_outs,
      outs_valid => buffer238_outs_valid,
      outs_ready => buffer238_outs_ready
    );

  addi17 : entity work.addi(arch) generic map(32)
    port map(
      lhs => buffer205_outs,
      lhs_valid => buffer205_outs_valid,
      lhs_ready => buffer205_outs_ready,
      rhs => buffer238_outs,
      rhs_valid => buffer238_outs_valid,
      rhs_ready => buffer238_outs_ready,
      clk => clk,
      rst => rst,
      result => addi17_result,
      result_valid => addi17_result_valid,
      result_ready => addi17_result_ready
    );

  buffer205 : entity work.tfifo(arch) generic map(3, 32)
    port map(
      ins => fork85_outs_2,
      ins_valid => fork85_outs_2_valid,
      ins_ready => fork85_outs_2_ready,
      clk => clk,
      rst => rst,
      outs => buffer205_outs,
      outs_valid => buffer205_outs_valid,
      outs_ready => buffer205_outs_ready
    );

  buffer239 : entity work.oehb_dataless(arch)
    port map(
      ins_valid => store5_doneOut_valid,
      ins_ready => store5_doneOut_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer239_outs_valid,
      outs_ready => buffer239_outs_ready
    );

  buffer5 : entity work.tfifo_dataless(arch) generic map(1)
    port map(
      ins_valid => buffer239_outs_valid,
      ins_ready => buffer239_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer5_outs_valid,
      outs_ready => buffer5_outs_ready
    );

  gate7 : entity work.gate(arch) generic map(2, 32)
    port map(
      ins(0) => addi17_result,
      ins_valid(0) => addi17_result_valid,
      ins_valid(1) => fork75_outs_0_valid,
      ins_ready(0) => addi17_result_ready,
      ins_ready(1) => fork75_outs_0_ready,
      clk => clk,
      rst => rst,
      outs => gate7_outs,
      outs_valid => gate7_outs_valid,
      outs_ready => gate7_outs_ready
    );

  trunci27 : entity work.trunci(arch) generic map(32, 7)
    port map(
      ins => gate7_outs,
      ins_valid => gate7_outs_valid,
      ins_ready => gate7_outs_ready,
      clk => clk,
      rst => rst,
      outs => trunci27_outs,
      outs_valid => trunci27_outs_valid,
      outs_ready => trunci27_outs_ready
    );

  store5 : entity work.store(arch) generic map(32, 7)
    port map(
      addrIn => trunci27_outs,
      addrIn_valid => trunci27_outs_valid,
      addrIn_ready => trunci27_outs_ready,
      dataIn => addi2_result,
      dataIn_valid => addi2_result_valid,
      dataIn_ready => addi2_result_ready,
      doneFromMem_valid => mem_controller4_stDone_1_valid,
      doneFromMem_ready => mem_controller4_stDone_1_ready,
      clk => clk,
      rst => rst,
      addrOut => store5_addrOut,
      addrOut_valid => store5_addrOut_valid,
      addrOut_ready => store5_addrOut_ready,
      dataToMem => store5_dataToMem,
      dataToMem_valid => store5_dataToMem_valid,
      dataToMem_ready => store5_dataToMem_ready,
      doneOut_valid => store5_doneOut_valid,
      doneOut_ready => store5_doneOut_ready
    );

  addi24 : entity work.addi(arch) generic map(6)
    port map(
      lhs => extsi88_outs,
      lhs_valid => extsi88_outs_valid,
      lhs_ready => extsi88_outs_ready,
      rhs => extsi93_outs,
      rhs_valid => extsi93_outs_valid,
      rhs_ready => extsi93_outs_ready,
      clk => clk,
      rst => rst,
      result => addi24_result,
      result_valid => addi24_result_valid,
      result_ready => addi24_result_ready
    );

  fork91 : entity work.handshake_fork(arch) generic map(2, 6)
    port map(
      ins => addi24_result,
      ins_valid => addi24_result_valid,
      ins_ready => addi24_result_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork91_outs_0,
      outs(1) => fork91_outs_1,
      outs_valid(0) => fork91_outs_0_valid,
      outs_valid(1) => fork91_outs_1_valid,
      outs_ready(0) => fork91_outs_0_ready,
      outs_ready(1) => fork91_outs_1_ready
    );

  trunci28 : entity work.trunci(arch) generic map(6, 5)
    port map(
      ins => buffer206_outs,
      ins_valid => buffer206_outs_valid,
      ins_ready => buffer206_outs_ready,
      clk => clk,
      rst => rst,
      outs => trunci28_outs,
      outs_valid => trunci28_outs_valid,
      outs_ready => trunci28_outs_ready
    );

  buffer206 : entity work.tfifo(arch) generic map(1, 6)
    port map(
      ins => fork91_outs_0,
      ins_valid => fork91_outs_0_valid,
      ins_ready => fork91_outs_0_ready,
      clk => clk,
      rst => rst,
      outs => buffer206_outs,
      outs_valid => buffer206_outs_valid,
      outs_ready => buffer206_outs_ready
    );

  buffer241 : entity work.oehb(arch) generic map(6)
    port map(
      ins => buffer207_outs,
      ins_valid => buffer207_outs_valid,
      ins_ready => buffer207_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer241_outs,
      outs_valid => buffer241_outs_valid,
      outs_ready => buffer241_outs_ready
    );

  cmpi6 : entity work.handshake_cmpi_0(arch) generic map(6)
    port map(
      lhs => buffer241_outs,
      lhs_valid => buffer241_outs_valid,
      lhs_ready => buffer241_outs_ready,
      rhs => extsi92_outs,
      rhs_valid => extsi92_outs_valid,
      rhs_ready => extsi92_outs_ready,
      clk => clk,
      rst => rst,
      result => cmpi6_result,
      result_valid => cmpi6_result_valid,
      result_ready => cmpi6_result_ready
    );

  buffer207 : entity work.tfifo(arch) generic map(1, 6)
    port map(
      ins => fork91_outs_1,
      ins_valid => fork91_outs_1_valid,
      ins_ready => fork91_outs_1_ready,
      clk => clk,
      rst => rst,
      outs => buffer207_outs,
      outs_valid => buffer207_outs_valid,
      outs_ready => buffer207_outs_ready
    );

  buffer240 : entity work.oehb(arch) generic map(1)
    port map(
      ins => cmpi6_result,
      ins_valid => cmpi6_result_valid,
      ins_ready => cmpi6_result_ready,
      clk => clk,
      rst => rst,
      outs => buffer240_outs,
      outs_valid => buffer240_outs_valid,
      outs_ready => buffer240_outs_ready
    );

  fork92 : entity work.handshake_fork(arch) generic map(11, 1)
    port map(
      ins => buffer240_outs,
      ins_valid => buffer240_outs_valid,
      ins_ready => buffer240_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork92_outs_0,
      outs(1) => fork92_outs_1,
      outs(2) => fork92_outs_2,
      outs(3) => fork92_outs_3,
      outs(4) => fork92_outs_4,
      outs(5) => fork92_outs_5,
      outs(6) => fork92_outs_6,
      outs(7) => fork92_outs_7,
      outs(8) => fork92_outs_8,
      outs(9) => fork92_outs_9,
      outs(10) => fork92_outs_10,
      outs_valid(0) => fork92_outs_0_valid,
      outs_valid(1) => fork92_outs_1_valid,
      outs_valid(2) => fork92_outs_2_valid,
      outs_valid(3) => fork92_outs_3_valid,
      outs_valid(4) => fork92_outs_4_valid,
      outs_valid(5) => fork92_outs_5_valid,
      outs_valid(6) => fork92_outs_6_valid,
      outs_valid(7) => fork92_outs_7_valid,
      outs_valid(8) => fork92_outs_8_valid,
      outs_valid(9) => fork92_outs_9_valid,
      outs_valid(10) => fork92_outs_10_valid,
      outs_ready(0) => fork92_outs_0_ready,
      outs_ready(1) => fork92_outs_1_ready,
      outs_ready(2) => fork92_outs_2_ready,
      outs_ready(3) => fork92_outs_3_ready,
      outs_ready(4) => fork92_outs_4_ready,
      outs_ready(5) => fork92_outs_5_ready,
      outs_ready(6) => fork92_outs_6_ready,
      outs_ready(7) => fork92_outs_7_ready,
      outs_ready(8) => fork92_outs_8_ready,
      outs_ready(9) => fork92_outs_9_ready,
      outs_ready(10) => fork92_outs_10_ready
    );

  cond_br29 : entity work.cond_br(arch) generic map(5)
    port map(
      condition => fork92_outs_0,
      condition_valid => fork92_outs_0_valid,
      condition_ready => fork92_outs_0_ready,
      data => trunci28_outs,
      data_valid => trunci28_outs_valid,
      data_ready => trunci28_outs_ready,
      clk => clk,
      rst => rst,
      trueOut => cond_br29_trueOut,
      trueOut_valid => cond_br29_trueOut_valid,
      trueOut_ready => cond_br29_trueOut_ready,
      falseOut => cond_br29_falseOut,
      falseOut_valid => cond_br29_falseOut_valid,
      falseOut_ready => cond_br29_falseOut_ready
    );

  sink23 : entity work.sink(arch) generic map(5)
    port map(
      ins => cond_br29_falseOut,
      ins_valid => cond_br29_falseOut_valid,
      ins_ready => cond_br29_falseOut_ready,
      clk => clk,
      rst => rst
    );

  cond_br30 : entity work.cond_br(arch) generic map(5)
    port map(
      condition => buffer209_outs,
      condition_valid => buffer209_outs_valid,
      condition_ready => buffer209_outs_ready,
      data => buffer210_outs,
      data_valid => buffer210_outs_valid,
      data_ready => buffer210_outs_ready,
      clk => clk,
      rst => rst,
      trueOut => cond_br30_trueOut,
      trueOut_valid => cond_br30_trueOut_valid,
      trueOut_ready => cond_br30_trueOut_ready,
      falseOut => cond_br30_falseOut,
      falseOut_valid => cond_br30_falseOut_valid,
      falseOut_ready => cond_br30_falseOut_ready
    );

  buffer209 : entity work.tfifo(arch) generic map(1, 1)
    port map(
      ins => fork92_outs_1,
      ins_valid => fork92_outs_1_valid,
      ins_ready => fork92_outs_1_ready,
      clk => clk,
      rst => rst,
      outs => buffer209_outs,
      outs_valid => buffer209_outs_valid,
      outs_ready => buffer209_outs_ready
    );

  buffer210 : entity work.tfifo(arch) generic map(1, 5)
    port map(
      ins => fork82_outs_0,
      ins_valid => fork82_outs_0_valid,
      ins_ready => fork82_outs_0_ready,
      clk => clk,
      rst => rst,
      outs => buffer210_outs,
      outs_valid => buffer210_outs_valid,
      outs_ready => buffer210_outs_ready
    );

  cond_br31 : entity work.cond_br(arch) generic map(5)
    port map(
      condition => fork92_outs_2,
      condition_valid => fork92_outs_2_valid,
      condition_ready => fork92_outs_2_ready,
      data => buffer212_outs,
      data_valid => buffer212_outs_valid,
      data_ready => buffer212_outs_ready,
      clk => clk,
      rst => rst,
      trueOut => cond_br31_trueOut,
      trueOut_valid => cond_br31_trueOut_valid,
      trueOut_ready => cond_br31_trueOut_ready,
      falseOut => cond_br31_falseOut,
      falseOut_valid => cond_br31_falseOut_valid,
      falseOut_ready => cond_br31_falseOut_ready
    );

  buffer212 : entity work.tfifo(arch) generic map(1, 5)
    port map(
      ins => fork84_outs_0,
      ins_valid => fork84_outs_0_valid,
      ins_ready => fork84_outs_0_ready,
      clk => clk,
      rst => rst,
      outs => buffer212_outs,
      outs_valid => buffer212_outs_valid,
      outs_ready => buffer212_outs_ready
    );

  cond_br32 : entity work.cond_br_dataless(arch)
    port map(
      condition => buffer213_outs,
      condition_valid => buffer213_outs_valid,
      condition_ready => buffer213_outs_ready,
      data_valid => fork87_outs_1_valid,
      data_ready => fork87_outs_1_ready,
      clk => clk,
      rst => rst,
      trueOut_valid => cond_br32_trueOut_valid,
      trueOut_ready => cond_br32_trueOut_ready,
      falseOut_valid => cond_br32_falseOut_valid,
      falseOut_ready => cond_br32_falseOut_ready
    );

  buffer213 : entity work.tfifo(arch) generic map(1, 1)
    port map(
      ins => fork92_outs_10,
      ins_valid => fork92_outs_10_valid,
      ins_ready => fork92_outs_10_ready,
      clk => clk,
      rst => rst,
      outs => buffer213_outs,
      outs_valid => buffer213_outs_valid,
      outs_ready => buffer213_outs_ready
    );

  cond_br134 : entity work.cond_br_dataless(arch)
    port map(
      condition => buffer214_outs,
      condition_valid => buffer214_outs_valid,
      condition_ready => buffer214_outs_ready,
      data_valid => cond_br132_falseOut_valid,
      data_ready => cond_br132_falseOut_ready,
      clk => clk,
      rst => rst,
      trueOut_valid => cond_br134_trueOut_valid,
      trueOut_ready => cond_br134_trueOut_ready,
      falseOut_valid => cond_br134_falseOut_valid,
      falseOut_ready => cond_br134_falseOut_ready
    );

  buffer214 : entity work.tfifo(arch) generic map(1, 1)
    port map(
      ins => fork94_outs_6,
      ins_valid => fork94_outs_6_valid,
      ins_ready => fork94_outs_6_ready,
      clk => clk,
      rst => rst,
      outs => buffer214_outs,
      outs_valid => buffer214_outs_valid,
      outs_ready => buffer214_outs_ready
    );

  cond_br135 : entity work.cond_br_dataless(arch)
    port map(
      condition => fork94_outs_5,
      condition_valid => fork94_outs_5_valid,
      condition_ready => fork94_outs_5_ready,
      data_valid => fork64_outs_0_valid,
      data_ready => fork64_outs_0_ready,
      clk => clk,
      rst => rst,
      trueOut_valid => cond_br135_trueOut_valid,
      trueOut_ready => cond_br135_trueOut_ready,
      falseOut_valid => cond_br135_falseOut_valid,
      falseOut_ready => cond_br135_falseOut_ready
    );

  sink24 : entity work.sink_dataless(arch)
    port map(
      ins_valid => cond_br135_falseOut_valid,
      ins_ready => cond_br135_falseOut_ready,
      clk => clk,
      rst => rst
    );

  cond_br136 : entity work.cond_br_dataless(arch)
    port map(
      condition => fork94_outs_4,
      condition_valid => fork94_outs_4_valid,
      condition_ready => fork94_outs_4_ready,
      data_valid => fork67_outs_0_valid,
      data_ready => fork67_outs_0_ready,
      clk => clk,
      rst => rst,
      trueOut_valid => cond_br136_trueOut_valid,
      trueOut_ready => cond_br136_trueOut_ready,
      falseOut_valid => cond_br136_falseOut_valid,
      falseOut_ready => cond_br136_falseOut_ready
    );

  sink25 : entity work.sink_dataless(arch)
    port map(
      ins_valid => cond_br136_falseOut_valid,
      ins_ready => cond_br136_falseOut_ready,
      clk => clk,
      rst => rst
    );

  cond_br137 : entity work.cond_br_dataless(arch)
    port map(
      condition => buffer217_outs,
      condition_valid => buffer217_outs_valid,
      condition_ready => buffer217_outs_ready,
      data_valid => fork65_outs_0_valid,
      data_ready => fork65_outs_0_ready,
      clk => clk,
      rst => rst,
      trueOut_valid => cond_br137_trueOut_valid,
      trueOut_ready => cond_br137_trueOut_ready,
      falseOut_valid => cond_br137_falseOut_valid,
      falseOut_ready => cond_br137_falseOut_ready
    );

  buffer217 : entity work.tfifo(arch) generic map(1, 1)
    port map(
      ins => fork94_outs_3,
      ins_valid => fork94_outs_3_valid,
      ins_ready => fork94_outs_3_ready,
      clk => clk,
      rst => rst,
      outs => buffer217_outs,
      outs_valid => buffer217_outs_valid,
      outs_ready => buffer217_outs_ready
    );

  sink26 : entity work.sink_dataless(arch)
    port map(
      ins_valid => cond_br137_falseOut_valid,
      ins_ready => cond_br137_falseOut_ready,
      clk => clk,
      rst => rst
    );

  cond_br138 : entity work.cond_br_dataless(arch)
    port map(
      condition => fork94_outs_2,
      condition_valid => fork94_outs_2_valid,
      condition_ready => fork94_outs_2_ready,
      data_valid => fork66_outs_0_valid,
      data_ready => fork66_outs_0_ready,
      clk => clk,
      rst => rst,
      trueOut_valid => cond_br138_trueOut_valid,
      trueOut_ready => cond_br138_trueOut_ready,
      falseOut_valid => cond_br138_falseOut_valid,
      falseOut_ready => cond_br138_falseOut_ready
    );

  sink27 : entity work.sink_dataless(arch)
    port map(
      ins_valid => cond_br138_falseOut_valid,
      ins_ready => cond_br138_falseOut_ready,
      clk => clk,
      rst => rst
    );

  extsi94 : entity work.extsi(arch) generic map(5, 6)
    port map(
      ins => cond_br31_falseOut,
      ins_valid => cond_br31_falseOut_valid,
      ins_ready => cond_br31_falseOut_ready,
      clk => clk,
      rst => rst,
      outs => extsi94_outs,
      outs_valid => extsi94_outs_valid,
      outs_ready => extsi94_outs_ready
    );

  source23 : entity work.source(arch)
    port map(
      clk => clk,
      rst => rst,
      outs_valid => source23_outs_valid,
      outs_ready => source23_outs_ready
    );

  constant83 : entity work.handshake_constant_3(arch) generic map(5)
    port map(
      ctrl_valid => source23_outs_valid,
      ctrl_ready => source23_outs_ready,
      clk => clk,
      rst => rst,
      outs => constant83_outs,
      outs_valid => constant83_outs_valid,
      outs_ready => constant83_outs_ready
    );

  extsi95 : entity work.extsi(arch) generic map(5, 6)
    port map(
      ins => constant83_outs,
      ins_valid => constant83_outs_valid,
      ins_ready => constant83_outs_ready,
      clk => clk,
      rst => rst,
      outs => extsi95_outs,
      outs_valid => extsi95_outs_valid,
      outs_ready => extsi95_outs_ready
    );

  source24 : entity work.source(arch)
    port map(
      clk => clk,
      rst => rst,
      outs_valid => source24_outs_valid,
      outs_ready => source24_outs_ready
    );

  constant84 : entity work.handshake_constant_1(arch) generic map(2)
    port map(
      ctrl_valid => source24_outs_valid,
      ctrl_ready => source24_outs_ready,
      clk => clk,
      rst => rst,
      outs => constant84_outs,
      outs_valid => constant84_outs_valid,
      outs_ready => constant84_outs_ready
    );

  extsi96 : entity work.extsi(arch) generic map(2, 6)
    port map(
      ins => constant84_outs,
      ins_valid => constant84_outs_valid,
      ins_ready => constant84_outs_ready,
      clk => clk,
      rst => rst,
      outs => extsi96_outs,
      outs_valid => extsi96_outs_valid,
      outs_ready => extsi96_outs_ready
    );

  addi25 : entity work.addi(arch) generic map(6)
    port map(
      lhs => extsi94_outs,
      lhs_valid => extsi94_outs_valid,
      lhs_ready => extsi94_outs_ready,
      rhs => extsi96_outs,
      rhs_valid => extsi96_outs_valid,
      rhs_ready => extsi96_outs_ready,
      clk => clk,
      rst => rst,
      result => addi25_result,
      result_valid => addi25_result_valid,
      result_ready => addi25_result_ready
    );

  buffer243 : entity work.oehb(arch) generic map(6)
    port map(
      ins => addi25_result,
      ins_valid => addi25_result_valid,
      ins_ready => addi25_result_ready,
      clk => clk,
      rst => rst,
      outs => buffer243_outs,
      outs_valid => buffer243_outs_valid,
      outs_ready => buffer243_outs_ready
    );

  fork93 : entity work.handshake_fork(arch) generic map(2, 6)
    port map(
      ins => buffer243_outs,
      ins_valid => buffer243_outs_valid,
      ins_ready => buffer243_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork93_outs_0,
      outs(1) => fork93_outs_1,
      outs_valid(0) => fork93_outs_0_valid,
      outs_valid(1) => fork93_outs_1_valid,
      outs_ready(0) => fork93_outs_0_ready,
      outs_ready(1) => fork93_outs_1_ready
    );

  trunci29 : entity work.trunci(arch) generic map(6, 5)
    port map(
      ins => buffer219_outs,
      ins_valid => buffer219_outs_valid,
      ins_ready => buffer219_outs_ready,
      clk => clk,
      rst => rst,
      outs => trunci29_outs,
      outs_valid => trunci29_outs_valid,
      outs_ready => trunci29_outs_ready
    );

  buffer219 : entity work.tfifo(arch) generic map(1, 6)
    port map(
      ins => fork93_outs_0,
      ins_valid => fork93_outs_0_valid,
      ins_ready => fork93_outs_0_ready,
      clk => clk,
      rst => rst,
      outs => buffer219_outs,
      outs_valid => buffer219_outs_valid,
      outs_ready => buffer219_outs_ready
    );

  cmpi7 : entity work.handshake_cmpi_0(arch) generic map(6)
    port map(
      lhs => fork93_outs_1,
      lhs_valid => fork93_outs_1_valid,
      lhs_ready => fork93_outs_1_ready,
      rhs => extsi95_outs,
      rhs_valid => extsi95_outs_valid,
      rhs_ready => extsi95_outs_ready,
      clk => clk,
      rst => rst,
      result => cmpi7_result,
      result_valid => cmpi7_result_valid,
      result_ready => cmpi7_result_ready
    );

  buffer244 : entity work.oehb(arch) generic map(1)
    port map(
      ins => cmpi7_result,
      ins_valid => cmpi7_result_valid,
      ins_ready => cmpi7_result_ready,
      clk => clk,
      rst => rst,
      outs => buffer244_outs,
      outs_valid => buffer244_outs_valid,
      outs_ready => buffer244_outs_ready
    );

  fork94 : entity work.handshake_fork(arch) generic map(9, 1)
    port map(
      ins => buffer244_outs,
      ins_valid => buffer244_outs_valid,
      ins_ready => buffer244_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork94_outs_0,
      outs(1) => fork94_outs_1,
      outs(2) => fork94_outs_2,
      outs(3) => fork94_outs_3,
      outs(4) => fork94_outs_4,
      outs(5) => fork94_outs_5,
      outs(6) => fork94_outs_6,
      outs(7) => fork94_outs_7,
      outs(8) => fork94_outs_8,
      outs_valid(0) => fork94_outs_0_valid,
      outs_valid(1) => fork94_outs_1_valid,
      outs_valid(2) => fork94_outs_2_valid,
      outs_valid(3) => fork94_outs_3_valid,
      outs_valid(4) => fork94_outs_4_valid,
      outs_valid(5) => fork94_outs_5_valid,
      outs_valid(6) => fork94_outs_6_valid,
      outs_valid(7) => fork94_outs_7_valid,
      outs_valid(8) => fork94_outs_8_valid,
      outs_ready(0) => fork94_outs_0_ready,
      outs_ready(1) => fork94_outs_1_ready,
      outs_ready(2) => fork94_outs_2_ready,
      outs_ready(3) => fork94_outs_3_ready,
      outs_ready(4) => fork94_outs_4_ready,
      outs_ready(5) => fork94_outs_5_ready,
      outs_ready(6) => fork94_outs_6_ready,
      outs_ready(7) => fork94_outs_7_ready,
      outs_ready(8) => fork94_outs_8_ready
    );

  cond_br33 : entity work.cond_br(arch) generic map(5)
    port map(
      condition => fork94_outs_0,
      condition_valid => fork94_outs_0_valid,
      condition_ready => fork94_outs_0_ready,
      data => trunci29_outs,
      data_valid => trunci29_outs_valid,
      data_ready => trunci29_outs_ready,
      clk => clk,
      rst => rst,
      trueOut => cond_br33_trueOut,
      trueOut_valid => cond_br33_trueOut_valid,
      trueOut_ready => cond_br33_trueOut_ready,
      falseOut => cond_br33_falseOut,
      falseOut_valid => cond_br33_falseOut_valid,
      falseOut_ready => cond_br33_falseOut_ready
    );

  sink29 : entity work.sink(arch) generic map(5)
    port map(
      ins => cond_br33_falseOut,
      ins_valid => cond_br33_falseOut_valid,
      ins_ready => cond_br33_falseOut_ready,
      clk => clk,
      rst => rst
    );

  cond_br34 : entity work.cond_br(arch) generic map(5)
    port map(
      condition => fork94_outs_1,
      condition_valid => fork94_outs_1_valid,
      condition_ready => fork94_outs_1_ready,
      data => cond_br30_falseOut,
      data_valid => cond_br30_falseOut_valid,
      data_ready => cond_br30_falseOut_ready,
      clk => clk,
      rst => rst,
      trueOut => cond_br34_trueOut,
      trueOut_valid => cond_br34_trueOut_valid,
      trueOut_ready => cond_br34_trueOut_ready,
      falseOut => cond_br34_falseOut,
      falseOut_valid => cond_br34_falseOut_valid,
      falseOut_ready => cond_br34_falseOut_ready
    );

  cond_br35 : entity work.cond_br_dataless(arch)
    port map(
      condition => buffer223_outs,
      condition_valid => buffer223_outs_valid,
      condition_ready => buffer223_outs_ready,
      data_valid => cond_br32_falseOut_valid,
      data_ready => cond_br32_falseOut_ready,
      clk => clk,
      rst => rst,
      trueOut_valid => cond_br35_trueOut_valid,
      trueOut_ready => cond_br35_trueOut_ready,
      falseOut_valid => cond_br35_falseOut_valid,
      falseOut_ready => cond_br35_falseOut_ready
    );

  buffer223 : entity work.tfifo(arch) generic map(1, 1)
    port map(
      ins => fork94_outs_8,
      ins_valid => fork94_outs_8_valid,
      ins_ready => fork94_outs_8_ready,
      clk => clk,
      rst => rst,
      outs => buffer223_outs,
      outs_valid => buffer223_outs_valid,
      outs_ready => buffer223_outs_ready
    );

  cond_br139 : entity work.cond_br_dataless(arch)
    port map(
      condition => fork96_outs_5,
      condition_valid => fork96_outs_5_valid,
      condition_ready => fork96_outs_5_ready,
      data_valid => fork58_outs_0_valid,
      data_ready => fork58_outs_0_ready,
      clk => clk,
      rst => rst,
      trueOut_valid => cond_br139_trueOut_valid,
      trueOut_ready => cond_br139_trueOut_ready,
      falseOut_valid => cond_br139_falseOut_valid,
      falseOut_ready => cond_br139_falseOut_ready
    );

  sink30 : entity work.sink_dataless(arch)
    port map(
      ins_valid => cond_br139_falseOut_valid,
      ins_ready => cond_br139_falseOut_ready,
      clk => clk,
      rst => rst
    );

  cond_br140 : entity work.cond_br_dataless(arch)
    port map(
      condition => buffer225_outs,
      condition_valid => buffer225_outs_valid,
      condition_ready => buffer225_outs_ready,
      data_valid => cond_br134_falseOut_valid,
      data_ready => cond_br134_falseOut_ready,
      clk => clk,
      rst => rst,
      trueOut_valid => cond_br140_trueOut_valid,
      trueOut_ready => cond_br140_trueOut_ready,
      falseOut_valid => cond_br140_falseOut_valid,
      falseOut_ready => cond_br140_falseOut_ready
    );

  buffer225 : entity work.tfifo(arch) generic map(1, 1)
    port map(
      ins => fork96_outs_4,
      ins_valid => fork96_outs_4_valid,
      ins_ready => fork96_outs_4_ready,
      clk => clk,
      rst => rst,
      outs => buffer225_outs,
      outs_valid => buffer225_outs_valid,
      outs_ready => buffer225_outs_ready
    );

  sink31 : entity work.sink_dataless(arch)
    port map(
      ins_valid => cond_br140_falseOut_valid,
      ins_ready => cond_br140_falseOut_ready,
      clk => clk,
      rst => rst
    );

  cond_br141 : entity work.cond_br_dataless(arch)
    port map(
      condition => fork96_outs_3,
      condition_valid => fork96_outs_3_valid,
      condition_ready => fork96_outs_3_ready,
      data_valid => fork60_outs_0_valid,
      data_ready => fork60_outs_0_ready,
      clk => clk,
      rst => rst,
      trueOut_valid => cond_br141_trueOut_valid,
      trueOut_ready => cond_br141_trueOut_ready,
      falseOut_valid => cond_br141_falseOut_valid,
      falseOut_ready => cond_br141_falseOut_ready
    );

  sink32 : entity work.sink_dataless(arch)
    port map(
      ins_valid => cond_br141_falseOut_valid,
      ins_ready => cond_br141_falseOut_ready,
      clk => clk,
      rst => rst
    );

  cond_br142 : entity work.cond_br_dataless(arch)
    port map(
      condition => fork96_outs_2,
      condition_valid => fork96_outs_2_valid,
      condition_ready => fork96_outs_2_ready,
      data_valid => fork59_outs_0_valid,
      data_ready => fork59_outs_0_ready,
      clk => clk,
      rst => rst,
      trueOut_valid => cond_br142_trueOut_valid,
      trueOut_ready => cond_br142_trueOut_ready,
      falseOut_valid => cond_br142_falseOut_valid,
      falseOut_ready => cond_br142_falseOut_ready
    );

  sink33 : entity work.sink_dataless(arch)
    port map(
      ins_valid => cond_br142_falseOut_valid,
      ins_ready => cond_br142_falseOut_ready,
      clk => clk,
      rst => rst
    );

  cond_br143 : entity work.cond_br_dataless(arch)
    port map(
      condition => fork96_outs_1,
      condition_valid => fork96_outs_1_valid,
      condition_ready => fork96_outs_1_ready,
      data_valid => fork61_outs_0_valid,
      data_ready => fork61_outs_0_ready,
      clk => clk,
      rst => rst,
      trueOut_valid => cond_br143_trueOut_valid,
      trueOut_ready => cond_br143_trueOut_ready,
      falseOut_valid => cond_br143_falseOut_valid,
      falseOut_ready => cond_br143_falseOut_ready
    );

  sink34 : entity work.sink_dataless(arch)
    port map(
      ins_valid => cond_br143_falseOut_valid,
      ins_ready => cond_br143_falseOut_ready,
      clk => clk,
      rst => rst
    );

  buffer246 : entity work.oehb(arch) generic map(5)
    port map(
      ins => cond_br34_falseOut,
      ins_valid => cond_br34_falseOut_valid,
      ins_ready => cond_br34_falseOut_ready,
      clk => clk,
      rst => rst,
      outs => buffer246_outs,
      outs_valid => buffer246_outs_valid,
      outs_ready => buffer246_outs_ready
    );

  extsi97 : entity work.extsi(arch) generic map(5, 6)
    port map(
      ins => buffer246_outs,
      ins_valid => buffer246_outs_valid,
      ins_ready => buffer246_outs_ready,
      clk => clk,
      rst => rst,
      outs => extsi97_outs,
      outs_valid => extsi97_outs_valid,
      outs_ready => extsi97_outs_ready
    );

  source25 : entity work.source(arch)
    port map(
      clk => clk,
      rst => rst,
      outs_valid => source25_outs_valid,
      outs_ready => source25_outs_ready
    );

  constant85 : entity work.handshake_constant_3(arch) generic map(5)
    port map(
      ctrl_valid => source25_outs_valid,
      ctrl_ready => source25_outs_ready,
      clk => clk,
      rst => rst,
      outs => constant85_outs,
      outs_valid => constant85_outs_valid,
      outs_ready => constant85_outs_ready
    );

  extsi98 : entity work.extsi(arch) generic map(5, 6)
    port map(
      ins => constant85_outs,
      ins_valid => constant85_outs_valid,
      ins_ready => constant85_outs_ready,
      clk => clk,
      rst => rst,
      outs => extsi98_outs,
      outs_valid => extsi98_outs_valid,
      outs_ready => extsi98_outs_ready
    );

  source26 : entity work.source(arch)
    port map(
      clk => clk,
      rst => rst,
      outs_valid => source26_outs_valid,
      outs_ready => source26_outs_ready
    );

  constant86 : entity work.handshake_constant_1(arch) generic map(2)
    port map(
      ctrl_valid => source26_outs_valid,
      ctrl_ready => source26_outs_ready,
      clk => clk,
      rst => rst,
      outs => constant86_outs,
      outs_valid => constant86_outs_valid,
      outs_ready => constant86_outs_ready
    );

  extsi99 : entity work.extsi(arch) generic map(2, 6)
    port map(
      ins => constant86_outs,
      ins_valid => constant86_outs_valid,
      ins_ready => constant86_outs_ready,
      clk => clk,
      rst => rst,
      outs => extsi99_outs,
      outs_valid => extsi99_outs_valid,
      outs_ready => extsi99_outs_ready
    );

  addi26 : entity work.addi(arch) generic map(6)
    port map(
      lhs => extsi97_outs,
      lhs_valid => extsi97_outs_valid,
      lhs_ready => extsi97_outs_ready,
      rhs => extsi99_outs,
      rhs_valid => extsi99_outs_valid,
      rhs_ready => extsi99_outs_ready,
      clk => clk,
      rst => rst,
      result => addi26_result,
      result_valid => addi26_result_valid,
      result_ready => addi26_result_ready
    );

  buffer247 : entity work.oehb(arch) generic map(6)
    port map(
      ins => addi26_result,
      ins_valid => addi26_result_valid,
      ins_ready => addi26_result_ready,
      clk => clk,
      rst => rst,
      outs => buffer247_outs,
      outs_valid => buffer247_outs_valid,
      outs_ready => buffer247_outs_ready
    );

  fork95 : entity work.handshake_fork(arch) generic map(2, 6)
    port map(
      ins => buffer247_outs,
      ins_valid => buffer247_outs_valid,
      ins_ready => buffer247_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork95_outs_0,
      outs(1) => fork95_outs_1,
      outs_valid(0) => fork95_outs_0_valid,
      outs_valid(1) => fork95_outs_1_valid,
      outs_ready(0) => fork95_outs_0_ready,
      outs_ready(1) => fork95_outs_1_ready
    );

  trunci30 : entity work.trunci(arch) generic map(6, 5)
    port map(
      ins => fork95_outs_0,
      ins_valid => fork95_outs_0_valid,
      ins_ready => fork95_outs_0_ready,
      clk => clk,
      rst => rst,
      outs => trunci30_outs,
      outs_valid => trunci30_outs_valid,
      outs_ready => trunci30_outs_ready
    );

  cmpi8 : entity work.handshake_cmpi_0(arch) generic map(6)
    port map(
      lhs => fork95_outs_1,
      lhs_valid => fork95_outs_1_valid,
      lhs_ready => fork95_outs_1_ready,
      rhs => extsi98_outs,
      rhs_valid => extsi98_outs_valid,
      rhs_ready => extsi98_outs_ready,
      clk => clk,
      rst => rst,
      result => cmpi8_result,
      result_valid => cmpi8_result_valid,
      result_ready => cmpi8_result_ready
    );

  buffer248 : entity work.oehb(arch) generic map(1)
    port map(
      ins => cmpi8_result,
      ins_valid => cmpi8_result_valid,
      ins_ready => cmpi8_result_ready,
      clk => clk,
      rst => rst,
      outs => buffer248_outs,
      outs_valid => buffer248_outs_valid,
      outs_ready => buffer248_outs_ready
    );

  fork96 : entity work.handshake_fork(arch) generic map(8, 1)
    port map(
      ins => buffer248_outs,
      ins_valid => buffer248_outs_valid,
      ins_ready => buffer248_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork96_outs_0,
      outs(1) => fork96_outs_1,
      outs(2) => fork96_outs_2,
      outs(3) => fork96_outs_3,
      outs(4) => fork96_outs_4,
      outs(5) => fork96_outs_5,
      outs(6) => fork96_outs_6,
      outs(7) => fork96_outs_7,
      outs_valid(0) => fork96_outs_0_valid,
      outs_valid(1) => fork96_outs_1_valid,
      outs_valid(2) => fork96_outs_2_valid,
      outs_valid(3) => fork96_outs_3_valid,
      outs_valid(4) => fork96_outs_4_valid,
      outs_valid(5) => fork96_outs_5_valid,
      outs_valid(6) => fork96_outs_6_valid,
      outs_valid(7) => fork96_outs_7_valid,
      outs_ready(0) => fork96_outs_0_ready,
      outs_ready(1) => fork96_outs_1_ready,
      outs_ready(2) => fork96_outs_2_ready,
      outs_ready(3) => fork96_outs_3_ready,
      outs_ready(4) => fork96_outs_4_ready,
      outs_ready(5) => fork96_outs_5_ready,
      outs_ready(6) => fork96_outs_6_ready,
      outs_ready(7) => fork96_outs_7_ready
    );

  cond_br36 : entity work.cond_br(arch) generic map(5)
    port map(
      condition => fork96_outs_0,
      condition_valid => fork96_outs_0_valid,
      condition_ready => fork96_outs_0_ready,
      data => trunci30_outs,
      data_valid => trunci30_outs_valid,
      data_ready => trunci30_outs_ready,
      clk => clk,
      rst => rst,
      trueOut => cond_br36_trueOut,
      trueOut_valid => cond_br36_trueOut_valid,
      trueOut_ready => cond_br36_trueOut_ready,
      falseOut => cond_br36_falseOut,
      falseOut_valid => cond_br36_falseOut_valid,
      falseOut_ready => cond_br36_falseOut_ready
    );

  sink36 : entity work.sink(arch) generic map(5)
    port map(
      ins => cond_br36_falseOut,
      ins_valid => cond_br36_falseOut_valid,
      ins_ready => cond_br36_falseOut_ready,
      clk => clk,
      rst => rst
    );

  cond_br37 : entity work.cond_br_dataless(arch)
    port map(
      condition => buffer232_outs,
      condition_valid => buffer232_outs_valid,
      condition_ready => buffer232_outs_ready,
      data_valid => cond_br35_falseOut_valid,
      data_ready => cond_br35_falseOut_ready,
      clk => clk,
      rst => rst,
      trueOut_valid => cond_br37_trueOut_valid,
      trueOut_ready => cond_br37_trueOut_ready,
      falseOut_valid => cond_br37_falseOut_valid,
      falseOut_ready => cond_br37_falseOut_ready
    );

  buffer232 : entity work.tfifo(arch) generic map(1, 1)
    port map(
      ins => fork96_outs_7,
      ins_valid => fork96_outs_7_valid,
      ins_ready => fork96_outs_7_ready,
      clk => clk,
      rst => rst,
      outs => buffer232_outs,
      outs_valid => buffer232_outs_valid,
      outs_ready => buffer232_outs_ready
    );

  fork97 : entity work.fork_dataless(arch) generic map(7)
    port map(
      ins_valid => cond_br37_falseOut_valid,
      ins_ready => cond_br37_falseOut_ready,
      clk => clk,
      rst => rst,
      outs_valid(0) => fork97_outs_0_valid,
      outs_valid(1) => fork97_outs_1_valid,
      outs_valid(2) => fork97_outs_2_valid,
      outs_valid(3) => fork97_outs_3_valid,
      outs_valid(4) => fork97_outs_4_valid,
      outs_valid(5) => fork97_outs_5_valid,
      outs_valid(6) => fork97_outs_6_valid,
      outs_ready(0) => fork97_outs_0_ready,
      outs_ready(1) => fork97_outs_1_ready,
      outs_ready(2) => fork97_outs_2_ready,
      outs_ready(3) => fork97_outs_3_ready,
      outs_ready(4) => fork97_outs_4_ready,
      outs_ready(5) => fork97_outs_5_ready,
      outs_ready(6) => fork97_outs_6_ready
    );

end architecture;
