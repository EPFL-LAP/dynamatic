library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity kernel_2mm is
  port (
    alpha : in std_logic_vector(31 downto 0);
    alpha_valid : in std_logic;
    beta : in std_logic_vector(31 downto 0);
    beta_valid : in std_logic;
    tmp_loadData : in std_logic_vector(31 downto 0);
    A_loadData : in std_logic_vector(31 downto 0);
    B_loadData : in std_logic_vector(31 downto 0);
    C_loadData : in std_logic_vector(31 downto 0);
    D_loadData : in std_logic_vector(31 downto 0);
    tmp_start_valid : in std_logic;
    A_start_valid : in std_logic;
    B_start_valid : in std_logic;
    C_start_valid : in std_logic;
    D_start_valid : in std_logic;
    start_valid : in std_logic;
    clk : in std_logic;
    rst : in std_logic;
    tmp_end_ready : in std_logic;
    A_end_ready : in std_logic;
    B_end_ready : in std_logic;
    C_end_ready : in std_logic;
    D_end_ready : in std_logic;
    end_ready : in std_logic;
    alpha_ready : out std_logic;
    beta_ready : out std_logic;
    tmp_start_ready : out std_logic;
    A_start_ready : out std_logic;
    B_start_ready : out std_logic;
    C_start_ready : out std_logic;
    D_start_ready : out std_logic;
    start_ready : out std_logic;
    tmp_end_valid : out std_logic;
    A_end_valid : out std_logic;
    B_end_valid : out std_logic;
    C_end_valid : out std_logic;
    D_end_valid : out std_logic;
    end_valid : out std_logic;
    tmp_loadEn : out std_logic;
    tmp_loadAddr : out std_logic_vector(6 downto 0);
    tmp_storeEn : out std_logic;
    tmp_storeAddr : out std_logic_vector(6 downto 0);
    tmp_storeData : out std_logic_vector(31 downto 0);
    A_loadEn : out std_logic;
    A_loadAddr : out std_logic_vector(6 downto 0);
    A_storeEn : out std_logic;
    A_storeAddr : out std_logic_vector(6 downto 0);
    A_storeData : out std_logic_vector(31 downto 0);
    B_loadEn : out std_logic;
    B_loadAddr : out std_logic_vector(6 downto 0);
    B_storeEn : out std_logic;
    B_storeAddr : out std_logic_vector(6 downto 0);
    B_storeData : out std_logic_vector(31 downto 0);
    C_loadEn : out std_logic;
    C_loadAddr : out std_logic_vector(6 downto 0);
    C_storeEn : out std_logic;
    C_storeAddr : out std_logic_vector(6 downto 0);
    C_storeData : out std_logic_vector(31 downto 0);
    D_loadEn : out std_logic;
    D_loadAddr : out std_logic_vector(6 downto 0);
    D_storeEn : out std_logic;
    D_storeAddr : out std_logic_vector(6 downto 0);
    D_storeData : out std_logic_vector(31 downto 0)
  );
end entity;

architecture behavioral of kernel_2mm is

  signal fork0_outs_0_valid : std_logic;
  signal fork0_outs_0_ready : std_logic;
  signal fork0_outs_1_valid : std_logic;
  signal fork0_outs_1_ready : std_logic;
  signal fork0_outs_2_valid : std_logic;
  signal fork0_outs_2_ready : std_logic;
  signal fork0_outs_3_valid : std_logic;
  signal fork0_outs_3_ready : std_logic;
  signal fork0_outs_4_valid : std_logic;
  signal fork0_outs_4_ready : std_logic;
  signal mem_controller3_ldData_0 : std_logic_vector(31 downto 0);
  signal mem_controller3_ldData_0_valid : std_logic;
  signal mem_controller3_ldData_0_ready : std_logic;
  signal mem_controller3_stDone_0_valid : std_logic;
  signal mem_controller3_stDone_0_ready : std_logic;
  signal mem_controller3_ldData_1 : std_logic_vector(31 downto 0);
  signal mem_controller3_ldData_1_valid : std_logic;
  signal mem_controller3_ldData_1_ready : std_logic;
  signal mem_controller3_stDone_1_valid : std_logic;
  signal mem_controller3_stDone_1_ready : std_logic;
  signal mem_controller3_memEnd_valid : std_logic;
  signal mem_controller3_memEnd_ready : std_logic;
  signal mem_controller3_loadEn : std_logic;
  signal mem_controller3_loadAddr : std_logic_vector(6 downto 0);
  signal mem_controller3_storeEn : std_logic;
  signal mem_controller3_storeAddr : std_logic_vector(6 downto 0);
  signal mem_controller3_storeData : std_logic_vector(31 downto 0);
  signal mem_controller4_ldData_0 : std_logic_vector(31 downto 0);
  signal mem_controller4_ldData_0_valid : std_logic;
  signal mem_controller4_ldData_0_ready : std_logic;
  signal mem_controller4_memEnd_valid : std_logic;
  signal mem_controller4_memEnd_ready : std_logic;
  signal mem_controller4_loadEn : std_logic;
  signal mem_controller4_loadAddr : std_logic_vector(6 downto 0);
  signal mem_controller4_storeEn : std_logic;
  signal mem_controller4_storeAddr : std_logic_vector(6 downto 0);
  signal mem_controller4_storeData : std_logic_vector(31 downto 0);
  signal mem_controller5_ldData_0 : std_logic_vector(31 downto 0);
  signal mem_controller5_ldData_0_valid : std_logic;
  signal mem_controller5_ldData_0_ready : std_logic;
  signal mem_controller5_memEnd_valid : std_logic;
  signal mem_controller5_memEnd_ready : std_logic;
  signal mem_controller5_loadEn : std_logic;
  signal mem_controller5_loadAddr : std_logic_vector(6 downto 0);
  signal mem_controller5_storeEn : std_logic;
  signal mem_controller5_storeAddr : std_logic_vector(6 downto 0);
  signal mem_controller5_storeData : std_logic_vector(31 downto 0);
  signal mem_controller6_ldData_0 : std_logic_vector(31 downto 0);
  signal mem_controller6_ldData_0_valid : std_logic;
  signal mem_controller6_ldData_0_ready : std_logic;
  signal mem_controller6_memEnd_valid : std_logic;
  signal mem_controller6_memEnd_ready : std_logic;
  signal mem_controller6_loadEn : std_logic;
  signal mem_controller6_loadAddr : std_logic_vector(6 downto 0);
  signal mem_controller6_storeEn : std_logic;
  signal mem_controller6_storeAddr : std_logic_vector(6 downto 0);
  signal mem_controller6_storeData : std_logic_vector(31 downto 0);
  signal mem_controller7_stDone_0_valid : std_logic;
  signal mem_controller7_stDone_0_ready : std_logic;
  signal mem_controller7_ldData_0 : std_logic_vector(31 downto 0);
  signal mem_controller7_ldData_0_valid : std_logic;
  signal mem_controller7_ldData_0_ready : std_logic;
  signal mem_controller7_stDone_1_valid : std_logic;
  signal mem_controller7_stDone_1_ready : std_logic;
  signal mem_controller7_ldData_1 : std_logic_vector(31 downto 0);
  signal mem_controller7_ldData_1_valid : std_logic;
  signal mem_controller7_ldData_1_ready : std_logic;
  signal mem_controller7_memEnd_valid : std_logic;
  signal mem_controller7_memEnd_ready : std_logic;
  signal mem_controller7_loadEn : std_logic;
  signal mem_controller7_loadAddr : std_logic_vector(6 downto 0);
  signal mem_controller7_storeEn : std_logic;
  signal mem_controller7_storeAddr : std_logic_vector(6 downto 0);
  signal mem_controller7_storeData : std_logic_vector(31 downto 0);
  signal constant29_outs : std_logic_vector(0 downto 0);
  signal constant29_outs_valid : std_logic;
  signal constant29_outs_ready : std_logic;
  signal extsi34_outs : std_logic_vector(4 downto 0);
  signal extsi34_outs_valid : std_logic;
  signal extsi34_outs_ready : std_logic;
  signal mux25_outs_valid : std_logic;
  signal mux25_outs_ready : std_logic;
  signal init0_outs : std_logic_vector(0 downto 0);
  signal init0_outs_valid : std_logic;
  signal init0_outs_ready : std_logic;
  signal mux0_outs : std_logic_vector(4 downto 0);
  signal mux0_outs_valid : std_logic;
  signal mux0_outs_ready : std_logic;
  signal mux1_outs : std_logic_vector(31 downto 0);
  signal mux1_outs_valid : std_logic;
  signal mux1_outs_ready : std_logic;
  signal buffer7_outs : std_logic_vector(0 downto 0);
  signal buffer7_outs_valid : std_logic;
  signal buffer7_outs_ready : std_logic;
  signal mux2_outs : std_logic_vector(31 downto 0);
  signal mux2_outs_valid : std_logic;
  signal mux2_outs_ready : std_logic;
  signal buffer8_outs : std_logic_vector(0 downto 0);
  signal buffer8_outs_valid : std_logic;
  signal buffer8_outs_ready : std_logic;
  signal control_merge0_outs_valid : std_logic;
  signal control_merge0_outs_ready : std_logic;
  signal control_merge0_index : std_logic_vector(0 downto 0);
  signal control_merge0_index_valid : std_logic;
  signal control_merge0_index_ready : std_logic;
  signal fork1_outs_0 : std_logic_vector(0 downto 0);
  signal fork1_outs_0_valid : std_logic;
  signal fork1_outs_0_ready : std_logic;
  signal fork1_outs_1 : std_logic_vector(0 downto 0);
  signal fork1_outs_1_valid : std_logic;
  signal fork1_outs_1_ready : std_logic;
  signal fork1_outs_2 : std_logic_vector(0 downto 0);
  signal fork1_outs_2_valid : std_logic;
  signal fork1_outs_2_ready : std_logic;
  signal fork2_outs_0_valid : std_logic;
  signal fork2_outs_0_ready : std_logic;
  signal fork2_outs_1_valid : std_logic;
  signal fork2_outs_1_ready : std_logic;
  signal constant30_outs : std_logic_vector(0 downto 0);
  signal constant30_outs_valid : std_logic;
  signal constant30_outs_ready : std_logic;
  signal extsi33_outs : std_logic_vector(4 downto 0);
  signal extsi33_outs_valid : std_logic;
  signal extsi33_outs_ready : std_logic;
  signal buffer10_outs : std_logic_vector(31 downto 0);
  signal buffer10_outs_valid : std_logic;
  signal buffer10_outs_ready : std_logic;
  signal buffer11_outs : std_logic_vector(31 downto 0);
  signal buffer11_outs_valid : std_logic;
  signal buffer11_outs_ready : std_logic;
  signal buffer14_outs : std_logic_vector(31 downto 0);
  signal buffer14_outs_valid : std_logic;
  signal buffer14_outs_ready : std_logic;
  signal buffer6_outs : std_logic_vector(4 downto 0);
  signal buffer6_outs_valid : std_logic;
  signal buffer6_outs_ready : std_logic;
  signal buffer5_outs_valid : std_logic;
  signal buffer5_outs_ready : std_logic;
  signal mux30_outs_valid : std_logic;
  signal mux30_outs_ready : std_logic;
  signal init5_outs : std_logic_vector(0 downto 0);
  signal init5_outs_valid : std_logic;
  signal init5_outs_ready : std_logic;
  signal buffer9_outs : std_logic_vector(0 downto 0);
  signal buffer9_outs_valid : std_logic;
  signal buffer9_outs_ready : std_logic;
  signal mux3_outs : std_logic_vector(4 downto 0);
  signal mux3_outs_valid : std_logic;
  signal mux3_outs_ready : std_logic;
  signal buffer18_outs : std_logic_vector(4 downto 0);
  signal buffer18_outs_valid : std_logic;
  signal buffer18_outs_ready : std_logic;
  signal fork3_outs_0 : std_logic_vector(4 downto 0);
  signal fork3_outs_0_valid : std_logic;
  signal fork3_outs_0_ready : std_logic;
  signal fork3_outs_1 : std_logic_vector(4 downto 0);
  signal fork3_outs_1_valid : std_logic;
  signal fork3_outs_1_ready : std_logic;
  signal extsi35_outs : std_logic_vector(6 downto 0);
  signal extsi35_outs_valid : std_logic;
  signal extsi35_outs_ready : std_logic;
  signal buffer15_outs : std_logic_vector(31 downto 0);
  signal buffer15_outs_valid : std_logic;
  signal buffer15_outs_ready : std_logic;
  signal mux4_outs : std_logic_vector(31 downto 0);
  signal mux4_outs_valid : std_logic;
  signal mux4_outs_ready : std_logic;
  signal buffer12_outs : std_logic_vector(0 downto 0);
  signal buffer12_outs_valid : std_logic;
  signal buffer12_outs_ready : std_logic;
  signal mux5_outs : std_logic_vector(31 downto 0);
  signal mux5_outs_valid : std_logic;
  signal mux5_outs_ready : std_logic;
  signal buffer13_outs : std_logic_vector(0 downto 0);
  signal buffer13_outs_valid : std_logic;
  signal buffer13_outs_ready : std_logic;
  signal mux6_outs : std_logic_vector(4 downto 0);
  signal mux6_outs_valid : std_logic;
  signal mux6_outs_ready : std_logic;
  signal buffer21_outs : std_logic_vector(4 downto 0);
  signal buffer21_outs_valid : std_logic;
  signal buffer21_outs_ready : std_logic;
  signal buffer24_outs : std_logic_vector(4 downto 0);
  signal buffer24_outs_valid : std_logic;
  signal buffer24_outs_ready : std_logic;
  signal fork4_outs_0 : std_logic_vector(4 downto 0);
  signal fork4_outs_0_valid : std_logic;
  signal fork4_outs_0_ready : std_logic;
  signal fork4_outs_1 : std_logic_vector(4 downto 0);
  signal fork4_outs_1_valid : std_logic;
  signal fork4_outs_1_ready : std_logic;
  signal extsi36_outs : std_logic_vector(31 downto 0);
  signal extsi36_outs_valid : std_logic;
  signal extsi36_outs_ready : std_logic;
  signal fork5_outs_0 : std_logic_vector(31 downto 0);
  signal fork5_outs_0_valid : std_logic;
  signal fork5_outs_0_ready : std_logic;
  signal fork5_outs_1 : std_logic_vector(31 downto 0);
  signal fork5_outs_1_valid : std_logic;
  signal fork5_outs_1_ready : std_logic;
  signal control_merge1_outs_valid : std_logic;
  signal control_merge1_outs_ready : std_logic;
  signal control_merge1_index : std_logic_vector(0 downto 0);
  signal control_merge1_index_valid : std_logic;
  signal control_merge1_index_ready : std_logic;
  signal fork6_outs_0 : std_logic_vector(0 downto 0);
  signal fork6_outs_0_valid : std_logic;
  signal fork6_outs_0_ready : std_logic;
  signal fork6_outs_1 : std_logic_vector(0 downto 0);
  signal fork6_outs_1_valid : std_logic;
  signal fork6_outs_1_ready : std_logic;
  signal fork6_outs_2 : std_logic_vector(0 downto 0);
  signal fork6_outs_2_valid : std_logic;
  signal fork6_outs_2_ready : std_logic;
  signal fork6_outs_3 : std_logic_vector(0 downto 0);
  signal fork6_outs_3_valid : std_logic;
  signal fork6_outs_3_ready : std_logic;
  signal fork7_outs_0_valid : std_logic;
  signal fork7_outs_0_ready : std_logic;
  signal fork7_outs_1_valid : std_logic;
  signal fork7_outs_1_ready : std_logic;
  signal fork7_outs_2_valid : std_logic;
  signal fork7_outs_2_ready : std_logic;
  signal constant31_outs : std_logic_vector(1 downto 0);
  signal constant31_outs_valid : std_logic;
  signal constant31_outs_ready : std_logic;
  signal extsi2_outs : std_logic_vector(31 downto 0);
  signal extsi2_outs_valid : std_logic;
  signal extsi2_outs_ready : std_logic;
  signal constant32_outs : std_logic_vector(0 downto 0);
  signal constant32_outs_valid : std_logic;
  signal constant32_outs_ready : std_logic;
  signal fork8_outs_0 : std_logic_vector(0 downto 0);
  signal fork8_outs_0_valid : std_logic;
  signal fork8_outs_0_ready : std_logic;
  signal fork8_outs_1 : std_logic_vector(0 downto 0);
  signal fork8_outs_1_valid : std_logic;
  signal fork8_outs_1_ready : std_logic;
  signal extsi4_outs : std_logic_vector(31 downto 0);
  signal extsi4_outs_valid : std_logic;
  signal extsi4_outs_ready : std_logic;
  signal source0_outs_valid : std_logic;
  signal source0_outs_ready : std_logic;
  signal constant33_outs : std_logic_vector(1 downto 0);
  signal constant33_outs_valid : std_logic;
  signal constant33_outs_ready : std_logic;
  signal extsi5_outs : std_logic_vector(31 downto 0);
  signal extsi5_outs_valid : std_logic;
  signal extsi5_outs_ready : std_logic;
  signal source1_outs_valid : std_logic;
  signal source1_outs_ready : std_logic;
  signal constant34_outs : std_logic_vector(2 downto 0);
  signal constant34_outs_valid : std_logic;
  signal constant34_outs_ready : std_logic;
  signal extsi6_outs : std_logic_vector(31 downto 0);
  signal extsi6_outs_valid : std_logic;
  signal extsi6_outs_ready : std_logic;
  signal shli0_result : std_logic_vector(31 downto 0);
  signal shli0_result_valid : std_logic;
  signal shli0_result_ready : std_logic;
  signal buffer27_outs : std_logic_vector(31 downto 0);
  signal buffer27_outs_valid : std_logic;
  signal buffer27_outs_ready : std_logic;
  signal trunci0_outs : std_logic_vector(6 downto 0);
  signal trunci0_outs_valid : std_logic;
  signal trunci0_outs_ready : std_logic;
  signal shli1_result : std_logic_vector(31 downto 0);
  signal shli1_result_valid : std_logic;
  signal shli1_result_ready : std_logic;
  signal buffer29_outs : std_logic_vector(31 downto 0);
  signal buffer29_outs_valid : std_logic;
  signal buffer29_outs_ready : std_logic;
  signal trunci1_outs : std_logic_vector(6 downto 0);
  signal trunci1_outs_valid : std_logic;
  signal trunci1_outs_ready : std_logic;
  signal addi19_result : std_logic_vector(6 downto 0);
  signal addi19_result_valid : std_logic;
  signal addi19_result_ready : std_logic;
  signal buffer30_outs : std_logic_vector(6 downto 0);
  signal buffer30_outs_valid : std_logic;
  signal buffer30_outs_ready : std_logic;
  signal addi2_result : std_logic_vector(6 downto 0);
  signal addi2_result_valid : std_logic;
  signal addi2_result_ready : std_logic;
  signal buffer0_outs_valid : std_logic;
  signal buffer0_outs_ready : std_logic;
  signal fork9_outs_0_valid : std_logic;
  signal fork9_outs_0_ready : std_logic;
  signal fork9_outs_1_valid : std_logic;
  signal fork9_outs_1_ready : std_logic;
  signal buffer31_outs : std_logic_vector(6 downto 0);
  signal buffer31_outs_valid : std_logic;
  signal buffer31_outs_ready : std_logic;
  signal store0_addrOut : std_logic_vector(6 downto 0);
  signal store0_addrOut_valid : std_logic;
  signal store0_addrOut_ready : std_logic;
  signal store0_dataToMem : std_logic_vector(31 downto 0);
  signal store0_dataToMem_valid : std_logic;
  signal store0_dataToMem_ready : std_logic;
  signal store0_doneOut_valid : std_logic;
  signal store0_doneOut_ready : std_logic;
  signal extsi32_outs : std_logic_vector(4 downto 0);
  signal extsi32_outs_valid : std_logic;
  signal extsi32_outs_ready : std_logic;
  signal buffer19_outs : std_logic_vector(31 downto 0);
  signal buffer19_outs_valid : std_logic;
  signal buffer19_outs_ready : std_logic;
  signal buffer20_outs : std_logic_vector(31 downto 0);
  signal buffer20_outs_valid : std_logic;
  signal buffer20_outs_ready : std_logic;
  signal cond_br83_trueOut_valid : std_logic;
  signal cond_br83_trueOut_ready : std_logic;
  signal cond_br83_falseOut_valid : std_logic;
  signal cond_br83_falseOut_ready : std_logic;
  signal buffer22_outs : std_logic_vector(0 downto 0);
  signal buffer22_outs_valid : std_logic;
  signal buffer22_outs_ready : std_logic;
  signal buffer100_outs_valid : std_logic;
  signal buffer100_outs_ready : std_logic;
  signal cond_br84_trueOut_valid : std_logic;
  signal cond_br84_trueOut_ready : std_logic;
  signal cond_br84_falseOut_valid : std_logic;
  signal cond_br84_falseOut_ready : std_logic;
  signal buffer23_outs : std_logic_vector(0 downto 0);
  signal buffer23_outs_valid : std_logic;
  signal buffer23_outs_ready : std_logic;
  signal init10_outs : std_logic_vector(0 downto 0);
  signal init10_outs_valid : std_logic;
  signal init10_outs_ready : std_logic;
  signal fork10_outs_0 : std_logic_vector(0 downto 0);
  signal fork10_outs_0_valid : std_logic;
  signal fork10_outs_0_ready : std_logic;
  signal fork10_outs_1 : std_logic_vector(0 downto 0);
  signal fork10_outs_1_valid : std_logic;
  signal fork10_outs_1_ready : std_logic;
  signal mux31_outs_valid : std_logic;
  signal mux31_outs_ready : std_logic;
  signal buffer25_outs : std_logic_vector(0 downto 0);
  signal buffer25_outs_valid : std_logic;
  signal buffer25_outs_ready : std_logic;
  signal buffer32_outs_valid : std_logic;
  signal buffer32_outs_ready : std_logic;
  signal buffer33_outs_valid : std_logic;
  signal buffer33_outs_ready : std_logic;
  signal fork11_outs_0_valid : std_logic;
  signal fork11_outs_0_ready : std_logic;
  signal fork11_outs_1_valid : std_logic;
  signal fork11_outs_1_ready : std_logic;
  signal fork11_outs_2_valid : std_logic;
  signal fork11_outs_2_ready : std_logic;
  signal buffer16_outs_valid : std_logic;
  signal buffer16_outs_ready : std_logic;
  signal buffer17_outs_valid : std_logic;
  signal buffer17_outs_ready : std_logic;
  signal mux34_outs_valid : std_logic;
  signal mux34_outs_ready : std_logic;
  signal buffer26_outs : std_logic_vector(0 downto 0);
  signal buffer26_outs_valid : std_logic;
  signal buffer26_outs_ready : std_logic;
  signal mux7_outs : std_logic_vector(4 downto 0);
  signal mux7_outs_valid : std_logic;
  signal mux7_outs_ready : std_logic;
  signal buffer40_outs : std_logic_vector(4 downto 0);
  signal buffer40_outs_valid : std_logic;
  signal buffer40_outs_ready : std_logic;
  signal buffer42_outs : std_logic_vector(4 downto 0);
  signal buffer42_outs_valid : std_logic;
  signal buffer42_outs_ready : std_logic;
  signal fork12_outs_0 : std_logic_vector(4 downto 0);
  signal fork12_outs_0_valid : std_logic;
  signal fork12_outs_0_ready : std_logic;
  signal fork12_outs_1 : std_logic_vector(4 downto 0);
  signal fork12_outs_1_valid : std_logic;
  signal fork12_outs_1_ready : std_logic;
  signal fork12_outs_2 : std_logic_vector(4 downto 0);
  signal fork12_outs_2_valid : std_logic;
  signal fork12_outs_2_ready : std_logic;
  signal extsi37_outs : std_logic_vector(6 downto 0);
  signal extsi37_outs_valid : std_logic;
  signal extsi37_outs_ready : std_logic;
  signal buffer28_outs : std_logic_vector(4 downto 0);
  signal buffer28_outs_valid : std_logic;
  signal buffer28_outs_ready : std_logic;
  signal extsi38_outs : std_logic_vector(5 downto 0);
  signal extsi38_outs_valid : std_logic;
  signal extsi38_outs_ready : std_logic;
  signal extsi39_outs : std_logic_vector(31 downto 0);
  signal extsi39_outs_valid : std_logic;
  signal extsi39_outs_ready : std_logic;
  signal fork13_outs_0 : std_logic_vector(31 downto 0);
  signal fork13_outs_0_valid : std_logic;
  signal fork13_outs_0_ready : std_logic;
  signal fork13_outs_1 : std_logic_vector(31 downto 0);
  signal fork13_outs_1_valid : std_logic;
  signal fork13_outs_1_ready : std_logic;
  signal mux8_outs : std_logic_vector(31 downto 0);
  signal mux8_outs_valid : std_logic;
  signal mux8_outs_ready : std_logic;
  signal buffer45_outs : std_logic_vector(31 downto 0);
  signal buffer45_outs_valid : std_logic;
  signal buffer45_outs_ready : std_logic;
  signal buffer47_outs : std_logic_vector(31 downto 0);
  signal buffer47_outs_valid : std_logic;
  signal buffer47_outs_ready : std_logic;
  signal fork14_outs_0 : std_logic_vector(31 downto 0);
  signal fork14_outs_0_valid : std_logic;
  signal fork14_outs_0_ready : std_logic;
  signal fork14_outs_1 : std_logic_vector(31 downto 0);
  signal fork14_outs_1_valid : std_logic;
  signal fork14_outs_1_ready : std_logic;
  signal mux9_outs : std_logic_vector(31 downto 0);
  signal mux9_outs_valid : std_logic;
  signal mux9_outs_ready : std_logic;
  signal mux10_outs : std_logic_vector(4 downto 0);
  signal mux10_outs_valid : std_logic;
  signal mux10_outs_ready : std_logic;
  signal buffer72_outs : std_logic_vector(4 downto 0);
  signal buffer72_outs_valid : std_logic;
  signal buffer72_outs_ready : std_logic;
  signal buffer73_outs : std_logic_vector(4 downto 0);
  signal buffer73_outs_valid : std_logic;
  signal buffer73_outs_ready : std_logic;
  signal fork15_outs_0 : std_logic_vector(4 downto 0);
  signal fork15_outs_0_valid : std_logic;
  signal fork15_outs_0_ready : std_logic;
  signal fork15_outs_1 : std_logic_vector(4 downto 0);
  signal fork15_outs_1_valid : std_logic;
  signal fork15_outs_1_ready : std_logic;
  signal extsi40_outs : std_logic_vector(31 downto 0);
  signal extsi40_outs_valid : std_logic;
  signal extsi40_outs_ready : std_logic;
  signal buffer34_outs : std_logic_vector(4 downto 0);
  signal buffer34_outs_valid : std_logic;
  signal buffer34_outs_ready : std_logic;
  signal fork16_outs_0 : std_logic_vector(31 downto 0);
  signal fork16_outs_0_valid : std_logic;
  signal fork16_outs_0_ready : std_logic;
  signal fork16_outs_1 : std_logic_vector(31 downto 0);
  signal fork16_outs_1_valid : std_logic;
  signal fork16_outs_1_ready : std_logic;
  signal fork16_outs_2 : std_logic_vector(31 downto 0);
  signal fork16_outs_2_valid : std_logic;
  signal fork16_outs_2_ready : std_logic;
  signal fork16_outs_3 : std_logic_vector(31 downto 0);
  signal fork16_outs_3_valid : std_logic;
  signal fork16_outs_3_ready : std_logic;
  signal fork16_outs_4 : std_logic_vector(31 downto 0);
  signal fork16_outs_4_valid : std_logic;
  signal fork16_outs_4_ready : std_logic;
  signal fork16_outs_5 : std_logic_vector(31 downto 0);
  signal fork16_outs_5_valid : std_logic;
  signal fork16_outs_5_ready : std_logic;
  signal mux11_outs : std_logic_vector(4 downto 0);
  signal mux11_outs_valid : std_logic;
  signal mux11_outs_ready : std_logic;
  signal buffer35_outs : std_logic_vector(0 downto 0);
  signal buffer35_outs_valid : std_logic;
  signal buffer35_outs_ready : std_logic;
  signal buffer74_outs : std_logic_vector(4 downto 0);
  signal buffer74_outs_valid : std_logic;
  signal buffer74_outs_ready : std_logic;
  signal buffer77_outs : std_logic_vector(4 downto 0);
  signal buffer77_outs_valid : std_logic;
  signal buffer77_outs_ready : std_logic;
  signal fork17_outs_0 : std_logic_vector(4 downto 0);
  signal fork17_outs_0_valid : std_logic;
  signal fork17_outs_0_ready : std_logic;
  signal fork17_outs_1 : std_logic_vector(4 downto 0);
  signal fork17_outs_1_valid : std_logic;
  signal fork17_outs_1_ready : std_logic;
  signal fork17_outs_2 : std_logic_vector(4 downto 0);
  signal fork17_outs_2_valid : std_logic;
  signal fork17_outs_2_ready : std_logic;
  signal extsi41_outs : std_logic_vector(6 downto 0);
  signal extsi41_outs_valid : std_logic;
  signal extsi41_outs_ready : std_logic;
  signal buffer36_outs : std_logic_vector(4 downto 0);
  signal buffer36_outs_valid : std_logic;
  signal buffer36_outs_ready : std_logic;
  signal extsi42_outs : std_logic_vector(31 downto 0);
  signal extsi42_outs_valid : std_logic;
  signal extsi42_outs_ready : std_logic;
  signal fork18_outs_0 : std_logic_vector(31 downto 0);
  signal fork18_outs_0_valid : std_logic;
  signal fork18_outs_0_ready : std_logic;
  signal fork18_outs_1 : std_logic_vector(31 downto 0);
  signal fork18_outs_1_valid : std_logic;
  signal fork18_outs_1_ready : std_logic;
  signal control_merge2_outs_valid : std_logic;
  signal control_merge2_outs_ready : std_logic;
  signal control_merge2_index : std_logic_vector(0 downto 0);
  signal control_merge2_index_valid : std_logic;
  signal control_merge2_index_ready : std_logic;
  signal fork19_outs_0 : std_logic_vector(0 downto 0);
  signal fork19_outs_0_valid : std_logic;
  signal fork19_outs_0_ready : std_logic;
  signal fork19_outs_1 : std_logic_vector(0 downto 0);
  signal fork19_outs_1_valid : std_logic;
  signal fork19_outs_1_ready : std_logic;
  signal fork19_outs_2 : std_logic_vector(0 downto 0);
  signal fork19_outs_2_valid : std_logic;
  signal fork19_outs_2_ready : std_logic;
  signal fork19_outs_3 : std_logic_vector(0 downto 0);
  signal fork19_outs_3_valid : std_logic;
  signal fork19_outs_3_ready : std_logic;
  signal fork19_outs_4 : std_logic_vector(0 downto 0);
  signal fork19_outs_4_valid : std_logic;
  signal fork19_outs_4_ready : std_logic;
  signal fork20_outs_0_valid : std_logic;
  signal fork20_outs_0_ready : std_logic;
  signal fork20_outs_1_valid : std_logic;
  signal fork20_outs_1_ready : std_logic;
  signal constant35_outs : std_logic_vector(1 downto 0);
  signal constant35_outs_valid : std_logic;
  signal constant35_outs_ready : std_logic;
  signal extsi7_outs : std_logic_vector(31 downto 0);
  signal extsi7_outs_valid : std_logic;
  signal extsi7_outs_ready : std_logic;
  signal source2_outs_valid : std_logic;
  signal source2_outs_ready : std_logic;
  signal constant36_outs : std_logic_vector(4 downto 0);
  signal constant36_outs_valid : std_logic;
  signal constant36_outs_ready : std_logic;
  signal extsi43_outs : std_logic_vector(5 downto 0);
  signal extsi43_outs_valid : std_logic;
  signal extsi43_outs_ready : std_logic;
  signal source3_outs_valid : std_logic;
  signal source3_outs_ready : std_logic;
  signal constant37_outs : std_logic_vector(1 downto 0);
  signal constant37_outs_valid : std_logic;
  signal constant37_outs_ready : std_logic;
  signal fork21_outs_0 : std_logic_vector(1 downto 0);
  signal fork21_outs_0_valid : std_logic;
  signal fork21_outs_0_ready : std_logic;
  signal fork21_outs_1 : std_logic_vector(1 downto 0);
  signal fork21_outs_1_valid : std_logic;
  signal fork21_outs_1_ready : std_logic;
  signal extsi44_outs : std_logic_vector(5 downto 0);
  signal extsi44_outs_valid : std_logic;
  signal extsi44_outs_ready : std_logic;
  signal buffer38_outs : std_logic_vector(1 downto 0);
  signal buffer38_outs_valid : std_logic;
  signal buffer38_outs_ready : std_logic;
  signal extsi9_outs : std_logic_vector(31 downto 0);
  signal extsi9_outs_valid : std_logic;
  signal extsi9_outs_ready : std_logic;
  signal buffer39_outs : std_logic_vector(1 downto 0);
  signal buffer39_outs_valid : std_logic;
  signal buffer39_outs_ready : std_logic;
  signal fork22_outs_0 : std_logic_vector(31 downto 0);
  signal fork22_outs_0_valid : std_logic;
  signal fork22_outs_0_ready : std_logic;
  signal fork22_outs_1 : std_logic_vector(31 downto 0);
  signal fork22_outs_1_valid : std_logic;
  signal fork22_outs_1_ready : std_logic;
  signal fork22_outs_2 : std_logic_vector(31 downto 0);
  signal fork22_outs_2_valid : std_logic;
  signal fork22_outs_2_ready : std_logic;
  signal fork22_outs_3 : std_logic_vector(31 downto 0);
  signal fork22_outs_3_valid : std_logic;
  signal fork22_outs_3_ready : std_logic;
  signal source4_outs_valid : std_logic;
  signal source4_outs_ready : std_logic;
  signal constant38_outs : std_logic_vector(2 downto 0);
  signal constant38_outs_valid : std_logic;
  signal constant38_outs_ready : std_logic;
  signal extsi10_outs : std_logic_vector(31 downto 0);
  signal extsi10_outs_valid : std_logic;
  signal extsi10_outs_ready : std_logic;
  signal fork23_outs_0 : std_logic_vector(31 downto 0);
  signal fork23_outs_0_valid : std_logic;
  signal fork23_outs_0_ready : std_logic;
  signal fork23_outs_1 : std_logic_vector(31 downto 0);
  signal fork23_outs_1_valid : std_logic;
  signal fork23_outs_1_ready : std_logic;
  signal fork23_outs_2 : std_logic_vector(31 downto 0);
  signal fork23_outs_2_valid : std_logic;
  signal fork23_outs_2_ready : std_logic;
  signal fork23_outs_3 : std_logic_vector(31 downto 0);
  signal fork23_outs_3_valid : std_logic;
  signal fork23_outs_3_ready : std_logic;
  signal shli2_result : std_logic_vector(31 downto 0);
  signal shli2_result_valid : std_logic;
  signal shli2_result_ready : std_logic;
  signal buffer41_outs : std_logic_vector(31 downto 0);
  signal buffer41_outs_valid : std_logic;
  signal buffer41_outs_ready : std_logic;
  signal buffer81_outs : std_logic_vector(31 downto 0);
  signal buffer81_outs_valid : std_logic;
  signal buffer81_outs_ready : std_logic;
  signal trunci2_outs : std_logic_vector(6 downto 0);
  signal trunci2_outs_valid : std_logic;
  signal trunci2_outs_ready : std_logic;
  signal shli3_result : std_logic_vector(31 downto 0);
  signal shli3_result_valid : std_logic;
  signal shli3_result_ready : std_logic;
  signal buffer43_outs : std_logic_vector(31 downto 0);
  signal buffer43_outs_valid : std_logic;
  signal buffer43_outs_ready : std_logic;
  signal buffer82_outs : std_logic_vector(31 downto 0);
  signal buffer82_outs_valid : std_logic;
  signal buffer82_outs_ready : std_logic;
  signal trunci3_outs : std_logic_vector(6 downto 0);
  signal trunci3_outs_valid : std_logic;
  signal trunci3_outs_ready : std_logic;
  signal addi20_result : std_logic_vector(6 downto 0);
  signal addi20_result_valid : std_logic;
  signal addi20_result_ready : std_logic;
  signal buffer83_outs : std_logic_vector(6 downto 0);
  signal buffer83_outs_valid : std_logic;
  signal buffer83_outs_ready : std_logic;
  signal addi3_result : std_logic_vector(6 downto 0);
  signal addi3_result_valid : std_logic;
  signal addi3_result_ready : std_logic;
  signal load0_addrOut : std_logic_vector(6 downto 0);
  signal load0_addrOut_valid : std_logic;
  signal load0_addrOut_ready : std_logic;
  signal load0_dataOut : std_logic_vector(31 downto 0);
  signal load0_dataOut_valid : std_logic;
  signal load0_dataOut_ready : std_logic;
  signal muli0_result : std_logic_vector(31 downto 0);
  signal muli0_result_valid : std_logic;
  signal muli0_result_ready : std_logic;
  signal buffer44_outs : std_logic_vector(31 downto 0);
  signal buffer44_outs_valid : std_logic;
  signal buffer44_outs_ready : std_logic;
  signal shli4_result : std_logic_vector(31 downto 0);
  signal shli4_result_valid : std_logic;
  signal shli4_result_ready : std_logic;
  signal buffer46_outs : std_logic_vector(31 downto 0);
  signal buffer46_outs_valid : std_logic;
  signal buffer46_outs_ready : std_logic;
  signal buffer84_outs : std_logic_vector(31 downto 0);
  signal buffer84_outs_valid : std_logic;
  signal buffer84_outs_ready : std_logic;
  signal trunci4_outs : std_logic_vector(6 downto 0);
  signal trunci4_outs_valid : std_logic;
  signal trunci4_outs_ready : std_logic;
  signal shli5_result : std_logic_vector(31 downto 0);
  signal shli5_result_valid : std_logic;
  signal shli5_result_ready : std_logic;
  signal buffer48_outs : std_logic_vector(31 downto 0);
  signal buffer48_outs_valid : std_logic;
  signal buffer48_outs_ready : std_logic;
  signal buffer85_outs : std_logic_vector(31 downto 0);
  signal buffer85_outs_valid : std_logic;
  signal buffer85_outs_ready : std_logic;
  signal trunci5_outs : std_logic_vector(6 downto 0);
  signal trunci5_outs_valid : std_logic;
  signal trunci5_outs_ready : std_logic;
  signal addi21_result : std_logic_vector(6 downto 0);
  signal addi21_result_valid : std_logic;
  signal addi21_result_ready : std_logic;
  signal buffer86_outs : std_logic_vector(6 downto 0);
  signal buffer86_outs_valid : std_logic;
  signal buffer86_outs_ready : std_logic;
  signal addi4_result : std_logic_vector(6 downto 0);
  signal addi4_result_valid : std_logic;
  signal addi4_result_ready : std_logic;
  signal load1_addrOut : std_logic_vector(6 downto 0);
  signal load1_addrOut_valid : std_logic;
  signal load1_addrOut_ready : std_logic;
  signal load1_dataOut : std_logic_vector(31 downto 0);
  signal load1_dataOut_valid : std_logic;
  signal load1_dataOut_ready : std_logic;
  signal muli1_result : std_logic_vector(31 downto 0);
  signal muli1_result_valid : std_logic;
  signal muli1_result_ready : std_logic;
  signal shli6_result : std_logic_vector(31 downto 0);
  signal shli6_result_valid : std_logic;
  signal shli6_result_ready : std_logic;
  signal buffer49_outs : std_logic_vector(31 downto 0);
  signal buffer49_outs_valid : std_logic;
  signal buffer49_outs_ready : std_logic;
  signal buffer50_outs : std_logic_vector(31 downto 0);
  signal buffer50_outs_valid : std_logic;
  signal buffer50_outs_ready : std_logic;
  signal shli7_result : std_logic_vector(31 downto 0);
  signal shli7_result_valid : std_logic;
  signal shli7_result_ready : std_logic;
  signal buffer51_outs : std_logic_vector(31 downto 0);
  signal buffer51_outs_valid : std_logic;
  signal buffer51_outs_ready : std_logic;
  signal buffer52_outs : std_logic_vector(31 downto 0);
  signal buffer52_outs_valid : std_logic;
  signal buffer52_outs_ready : std_logic;
  signal buffer87_outs : std_logic_vector(31 downto 0);
  signal buffer87_outs_valid : std_logic;
  signal buffer87_outs_ready : std_logic;
  signal buffer88_outs : std_logic_vector(31 downto 0);
  signal buffer88_outs_valid : std_logic;
  signal buffer88_outs_ready : std_logic;
  signal addi22_result : std_logic_vector(31 downto 0);
  signal addi22_result_valid : std_logic;
  signal addi22_result_ready : std_logic;
  signal buffer92_outs : std_logic_vector(31 downto 0);
  signal buffer92_outs_valid : std_logic;
  signal buffer92_outs_ready : std_logic;
  signal addi5_result : std_logic_vector(31 downto 0);
  signal addi5_result_valid : std_logic;
  signal addi5_result_ready : std_logic;
  signal buffer53_outs : std_logic_vector(31 downto 0);
  signal buffer53_outs_valid : std_logic;
  signal buffer53_outs_ready : std_logic;
  signal buffer37_outs_valid : std_logic;
  signal buffer37_outs_ready : std_logic;
  signal gate0_outs : std_logic_vector(31 downto 0);
  signal gate0_outs_valid : std_logic;
  signal gate0_outs_ready : std_logic;
  signal trunci6_outs : std_logic_vector(6 downto 0);
  signal trunci6_outs_valid : std_logic;
  signal trunci6_outs_ready : std_logic;
  signal load2_addrOut : std_logic_vector(6 downto 0);
  signal load2_addrOut_valid : std_logic;
  signal load2_addrOut_ready : std_logic;
  signal load2_dataOut : std_logic_vector(31 downto 0);
  signal load2_dataOut_valid : std_logic;
  signal load2_dataOut_ready : std_logic;
  signal addi0_result : std_logic_vector(31 downto 0);
  signal addi0_result_valid : std_logic;
  signal addi0_result_ready : std_logic;
  signal shli8_result : std_logic_vector(31 downto 0);
  signal shli8_result_valid : std_logic;
  signal shli8_result_ready : std_logic;
  signal buffer54_outs : std_logic_vector(31 downto 0);
  signal buffer54_outs_valid : std_logic;
  signal buffer54_outs_ready : std_logic;
  signal buffer55_outs : std_logic_vector(31 downto 0);
  signal buffer55_outs_valid : std_logic;
  signal buffer55_outs_ready : std_logic;
  signal shli9_result : std_logic_vector(31 downto 0);
  signal shli9_result_valid : std_logic;
  signal shli9_result_ready : std_logic;
  signal buffer56_outs : std_logic_vector(31 downto 0);
  signal buffer56_outs_valid : std_logic;
  signal buffer56_outs_ready : std_logic;
  signal buffer57_outs : std_logic_vector(31 downto 0);
  signal buffer57_outs_valid : std_logic;
  signal buffer57_outs_ready : std_logic;
  signal buffer93_outs : std_logic_vector(31 downto 0);
  signal buffer93_outs_valid : std_logic;
  signal buffer93_outs_ready : std_logic;
  signal buffer94_outs : std_logic_vector(31 downto 0);
  signal buffer94_outs_valid : std_logic;
  signal buffer94_outs_ready : std_logic;
  signal addi23_result : std_logic_vector(31 downto 0);
  signal addi23_result_valid : std_logic;
  signal addi23_result_ready : std_logic;
  signal buffer99_outs : std_logic_vector(31 downto 0);
  signal buffer99_outs_valid : std_logic;
  signal buffer99_outs_ready : std_logic;
  signal addi6_result : std_logic_vector(31 downto 0);
  signal addi6_result_valid : std_logic;
  signal addi6_result_ready : std_logic;
  signal buffer58_outs : std_logic_vector(31 downto 0);
  signal buffer58_outs_valid : std_logic;
  signal buffer58_outs_ready : std_logic;
  signal buffer1_outs_valid : std_logic;
  signal buffer1_outs_ready : std_logic;
  signal gate1_outs : std_logic_vector(31 downto 0);
  signal gate1_outs_valid : std_logic;
  signal gate1_outs_ready : std_logic;
  signal trunci7_outs : std_logic_vector(6 downto 0);
  signal trunci7_outs_valid : std_logic;
  signal trunci7_outs_ready : std_logic;
  signal store1_addrOut : std_logic_vector(6 downto 0);
  signal store1_addrOut_valid : std_logic;
  signal store1_addrOut_ready : std_logic;
  signal store1_dataToMem : std_logic_vector(31 downto 0);
  signal store1_dataToMem_valid : std_logic;
  signal store1_dataToMem_ready : std_logic;
  signal store1_doneOut_valid : std_logic;
  signal store1_doneOut_ready : std_logic;
  signal addi13_result : std_logic_vector(5 downto 0);
  signal addi13_result_valid : std_logic;
  signal addi13_result_ready : std_logic;
  signal fork24_outs_0 : std_logic_vector(5 downto 0);
  signal fork24_outs_0_valid : std_logic;
  signal fork24_outs_0_ready : std_logic;
  signal fork24_outs_1 : std_logic_vector(5 downto 0);
  signal fork24_outs_1_valid : std_logic;
  signal fork24_outs_1_ready : std_logic;
  signal trunci8_outs : std_logic_vector(4 downto 0);
  signal trunci8_outs_valid : std_logic;
  signal trunci8_outs_ready : std_logic;
  signal buffer59_outs : std_logic_vector(5 downto 0);
  signal buffer59_outs_valid : std_logic;
  signal buffer59_outs_ready : std_logic;
  signal buffer103_outs : std_logic_vector(5 downto 0);
  signal buffer103_outs_valid : std_logic;
  signal buffer103_outs_ready : std_logic;
  signal cmpi0_result : std_logic_vector(0 downto 0);
  signal cmpi0_result_valid : std_logic;
  signal cmpi0_result_ready : std_logic;
  signal buffer60_outs : std_logic_vector(5 downto 0);
  signal buffer60_outs_valid : std_logic;
  signal buffer60_outs_ready : std_logic;
  signal buffer102_outs : std_logic_vector(0 downto 0);
  signal buffer102_outs_valid : std_logic;
  signal buffer102_outs_ready : std_logic;
  signal fork25_outs_0 : std_logic_vector(0 downto 0);
  signal fork25_outs_0_valid : std_logic;
  signal fork25_outs_0_ready : std_logic;
  signal fork25_outs_1 : std_logic_vector(0 downto 0);
  signal fork25_outs_1_valid : std_logic;
  signal fork25_outs_1_ready : std_logic;
  signal fork25_outs_2 : std_logic_vector(0 downto 0);
  signal fork25_outs_2_valid : std_logic;
  signal fork25_outs_2_ready : std_logic;
  signal fork25_outs_3 : std_logic_vector(0 downto 0);
  signal fork25_outs_3_valid : std_logic;
  signal fork25_outs_3_ready : std_logic;
  signal fork25_outs_4 : std_logic_vector(0 downto 0);
  signal fork25_outs_4_valid : std_logic;
  signal fork25_outs_4_ready : std_logic;
  signal fork25_outs_5 : std_logic_vector(0 downto 0);
  signal fork25_outs_5_valid : std_logic;
  signal fork25_outs_5_ready : std_logic;
  signal fork25_outs_6 : std_logic_vector(0 downto 0);
  signal fork25_outs_6_valid : std_logic;
  signal fork25_outs_6_ready : std_logic;
  signal fork25_outs_7 : std_logic_vector(0 downto 0);
  signal fork25_outs_7_valid : std_logic;
  signal fork25_outs_7_ready : std_logic;
  signal fork25_outs_8 : std_logic_vector(0 downto 0);
  signal fork25_outs_8_valid : std_logic;
  signal fork25_outs_8_ready : std_logic;
  signal cond_br6_trueOut : std_logic_vector(4 downto 0);
  signal cond_br6_trueOut_valid : std_logic;
  signal cond_br6_trueOut_ready : std_logic;
  signal cond_br6_falseOut : std_logic_vector(4 downto 0);
  signal cond_br6_falseOut_valid : std_logic;
  signal cond_br6_falseOut_ready : std_logic;
  signal cond_br7_trueOut : std_logic_vector(31 downto 0);
  signal cond_br7_trueOut_valid : std_logic;
  signal cond_br7_trueOut_ready : std_logic;
  signal cond_br7_falseOut : std_logic_vector(31 downto 0);
  signal cond_br7_falseOut_valid : std_logic;
  signal cond_br7_falseOut_ready : std_logic;
  signal buffer62_outs : std_logic_vector(0 downto 0);
  signal buffer62_outs_valid : std_logic;
  signal buffer62_outs_ready : std_logic;
  signal buffer63_outs : std_logic_vector(31 downto 0);
  signal buffer63_outs_valid : std_logic;
  signal buffer63_outs_ready : std_logic;
  signal buffer61_outs : std_logic_vector(31 downto 0);
  signal buffer61_outs_valid : std_logic;
  signal buffer61_outs_ready : std_logic;
  signal buffer67_outs : std_logic_vector(31 downto 0);
  signal buffer67_outs_valid : std_logic;
  signal buffer67_outs_ready : std_logic;
  signal cond_br8_trueOut : std_logic_vector(31 downto 0);
  signal cond_br8_trueOut_valid : std_logic;
  signal cond_br8_trueOut_ready : std_logic;
  signal cond_br8_falseOut : std_logic_vector(31 downto 0);
  signal cond_br8_falseOut_valid : std_logic;
  signal cond_br8_falseOut_ready : std_logic;
  signal buffer64_outs : std_logic_vector(0 downto 0);
  signal buffer64_outs_valid : std_logic;
  signal buffer64_outs_ready : std_logic;
  signal cond_br9_trueOut : std_logic_vector(4 downto 0);
  signal cond_br9_trueOut_valid : std_logic;
  signal cond_br9_trueOut_ready : std_logic;
  signal cond_br9_falseOut : std_logic_vector(4 downto 0);
  signal cond_br9_falseOut_valid : std_logic;
  signal cond_br9_falseOut_ready : std_logic;
  signal buffer65_outs : std_logic_vector(0 downto 0);
  signal buffer65_outs_valid : std_logic;
  signal buffer65_outs_ready : std_logic;
  signal buffer66_outs : std_logic_vector(4 downto 0);
  signal buffer66_outs_valid : std_logic;
  signal buffer66_outs_ready : std_logic;
  signal cond_br10_trueOut : std_logic_vector(4 downto 0);
  signal cond_br10_trueOut_valid : std_logic;
  signal cond_br10_trueOut_ready : std_logic;
  signal cond_br10_falseOut : std_logic_vector(4 downto 0);
  signal cond_br10_falseOut_valid : std_logic;
  signal cond_br10_falseOut_ready : std_logic;
  signal buffer68_outs : std_logic_vector(4 downto 0);
  signal buffer68_outs_valid : std_logic;
  signal buffer68_outs_ready : std_logic;
  signal buffer79_outs_valid : std_logic;
  signal buffer79_outs_ready : std_logic;
  signal cond_br11_trueOut_valid : std_logic;
  signal cond_br11_trueOut_ready : std_logic;
  signal cond_br11_falseOut_valid : std_logic;
  signal cond_br11_falseOut_ready : std_logic;
  signal buffer69_outs : std_logic_vector(0 downto 0);
  signal buffer69_outs_valid : std_logic;
  signal buffer69_outs_ready : std_logic;
  signal cond_br85_trueOut_valid : std_logic;
  signal cond_br85_trueOut_ready : std_logic;
  signal cond_br85_falseOut_valid : std_logic;
  signal cond_br85_falseOut_ready : std_logic;
  signal buffer70_outs : std_logic_vector(0 downto 0);
  signal buffer70_outs_valid : std_logic;
  signal buffer70_outs_ready : std_logic;
  signal cond_br86_trueOut_valid : std_logic;
  signal cond_br86_trueOut_ready : std_logic;
  signal cond_br86_falseOut_valid : std_logic;
  signal cond_br86_falseOut_ready : std_logic;
  signal buffer71_outs : std_logic_vector(0 downto 0);
  signal buffer71_outs_valid : std_logic;
  signal buffer71_outs_ready : std_logic;
  signal extsi45_outs : std_logic_vector(5 downto 0);
  signal extsi45_outs_valid : std_logic;
  signal extsi45_outs_ready : std_logic;
  signal source5_outs_valid : std_logic;
  signal source5_outs_ready : std_logic;
  signal constant39_outs : std_logic_vector(4 downto 0);
  signal constant39_outs_valid : std_logic;
  signal constant39_outs_ready : std_logic;
  signal extsi46_outs : std_logic_vector(5 downto 0);
  signal extsi46_outs_valid : std_logic;
  signal extsi46_outs_ready : std_logic;
  signal source6_outs_valid : std_logic;
  signal source6_outs_ready : std_logic;
  signal constant40_outs : std_logic_vector(1 downto 0);
  signal constant40_outs_valid : std_logic;
  signal constant40_outs_ready : std_logic;
  signal extsi47_outs : std_logic_vector(5 downto 0);
  signal extsi47_outs_valid : std_logic;
  signal extsi47_outs_ready : std_logic;
  signal addi14_result : std_logic_vector(5 downto 0);
  signal addi14_result_valid : std_logic;
  signal addi14_result_ready : std_logic;
  signal buffer106_outs : std_logic_vector(5 downto 0);
  signal buffer106_outs_valid : std_logic;
  signal buffer106_outs_ready : std_logic;
  signal fork26_outs_0 : std_logic_vector(5 downto 0);
  signal fork26_outs_0_valid : std_logic;
  signal fork26_outs_0_ready : std_logic;
  signal fork26_outs_1 : std_logic_vector(5 downto 0);
  signal fork26_outs_1_valid : std_logic;
  signal fork26_outs_1_ready : std_logic;
  signal trunci9_outs : std_logic_vector(4 downto 0);
  signal trunci9_outs_valid : std_logic;
  signal trunci9_outs_ready : std_logic;
  signal cmpi1_result : std_logic_vector(0 downto 0);
  signal cmpi1_result_valid : std_logic;
  signal cmpi1_result_ready : std_logic;
  signal buffer107_outs : std_logic_vector(0 downto 0);
  signal buffer107_outs_valid : std_logic;
  signal buffer107_outs_ready : std_logic;
  signal fork27_outs_0 : std_logic_vector(0 downto 0);
  signal fork27_outs_0_valid : std_logic;
  signal fork27_outs_0_ready : std_logic;
  signal fork27_outs_1 : std_logic_vector(0 downto 0);
  signal fork27_outs_1_valid : std_logic;
  signal fork27_outs_1_ready : std_logic;
  signal fork27_outs_2 : std_logic_vector(0 downto 0);
  signal fork27_outs_2_valid : std_logic;
  signal fork27_outs_2_ready : std_logic;
  signal fork27_outs_3 : std_logic_vector(0 downto 0);
  signal fork27_outs_3_valid : std_logic;
  signal fork27_outs_3_ready : std_logic;
  signal fork27_outs_4 : std_logic_vector(0 downto 0);
  signal fork27_outs_4_valid : std_logic;
  signal fork27_outs_4_ready : std_logic;
  signal fork27_outs_5 : std_logic_vector(0 downto 0);
  signal fork27_outs_5_valid : std_logic;
  signal fork27_outs_5_ready : std_logic;
  signal fork27_outs_6 : std_logic_vector(0 downto 0);
  signal fork27_outs_6_valid : std_logic;
  signal fork27_outs_6_ready : std_logic;
  signal fork27_outs_7 : std_logic_vector(0 downto 0);
  signal fork27_outs_7_valid : std_logic;
  signal fork27_outs_7_ready : std_logic;
  signal cond_br12_trueOut : std_logic_vector(4 downto 0);
  signal cond_br12_trueOut_valid : std_logic;
  signal cond_br12_trueOut_ready : std_logic;
  signal cond_br12_falseOut : std_logic_vector(4 downto 0);
  signal cond_br12_falseOut_valid : std_logic;
  signal cond_br12_falseOut_ready : std_logic;
  signal buffer104_outs : std_logic_vector(31 downto 0);
  signal buffer104_outs_valid : std_logic;
  signal buffer104_outs_ready : std_logic;
  signal cond_br13_trueOut : std_logic_vector(31 downto 0);
  signal cond_br13_trueOut_valid : std_logic;
  signal cond_br13_trueOut_ready : std_logic;
  signal cond_br13_falseOut : std_logic_vector(31 downto 0);
  signal cond_br13_falseOut_valid : std_logic;
  signal cond_br13_falseOut_ready : std_logic;
  signal buffer75_outs : std_logic_vector(0 downto 0);
  signal buffer75_outs_valid : std_logic;
  signal buffer75_outs_ready : std_logic;
  signal buffer105_outs : std_logic_vector(31 downto 0);
  signal buffer105_outs_valid : std_logic;
  signal buffer105_outs_ready : std_logic;
  signal cond_br14_trueOut : std_logic_vector(31 downto 0);
  signal cond_br14_trueOut_valid : std_logic;
  signal cond_br14_trueOut_ready : std_logic;
  signal cond_br14_falseOut : std_logic_vector(31 downto 0);
  signal cond_br14_falseOut_valid : std_logic;
  signal cond_br14_falseOut_ready : std_logic;
  signal buffer76_outs : std_logic_vector(0 downto 0);
  signal buffer76_outs_valid : std_logic;
  signal buffer76_outs_ready : std_logic;
  signal cond_br15_trueOut : std_logic_vector(4 downto 0);
  signal cond_br15_trueOut_valid : std_logic;
  signal cond_br15_trueOut_ready : std_logic;
  signal cond_br15_falseOut : std_logic_vector(4 downto 0);
  signal cond_br15_falseOut_valid : std_logic;
  signal cond_br15_falseOut_ready : std_logic;
  signal cond_br16_trueOut_valid : std_logic;
  signal cond_br16_trueOut_ready : std_logic;
  signal cond_br16_falseOut_valid : std_logic;
  signal cond_br16_falseOut_ready : std_logic;
  signal buffer78_outs : std_logic_vector(0 downto 0);
  signal buffer78_outs_valid : std_logic;
  signal buffer78_outs_ready : std_logic;
  signal cond_br87_trueOut_valid : std_logic;
  signal cond_br87_trueOut_ready : std_logic;
  signal cond_br87_falseOut_valid : std_logic;
  signal cond_br87_falseOut_ready : std_logic;
  signal cond_br88_trueOut_valid : std_logic;
  signal cond_br88_trueOut_ready : std_logic;
  signal cond_br88_falseOut_valid : std_logic;
  signal cond_br88_falseOut_ready : std_logic;
  signal buffer80_outs : std_logic_vector(0 downto 0);
  signal buffer80_outs_valid : std_logic;
  signal buffer80_outs_ready : std_logic;
  signal buffer108_outs : std_logic_vector(4 downto 0);
  signal buffer108_outs_valid : std_logic;
  signal buffer108_outs_ready : std_logic;
  signal extsi48_outs : std_logic_vector(5 downto 0);
  signal extsi48_outs_valid : std_logic;
  signal extsi48_outs_ready : std_logic;
  signal fork28_outs_0_valid : std_logic;
  signal fork28_outs_0_ready : std_logic;
  signal fork28_outs_1_valid : std_logic;
  signal fork28_outs_1_ready : std_logic;
  signal constant41_outs : std_logic_vector(0 downto 0);
  signal constant41_outs_valid : std_logic;
  signal constant41_outs_ready : std_logic;
  signal source7_outs_valid : std_logic;
  signal source7_outs_ready : std_logic;
  signal constant42_outs : std_logic_vector(4 downto 0);
  signal constant42_outs_valid : std_logic;
  signal constant42_outs_ready : std_logic;
  signal extsi49_outs : std_logic_vector(5 downto 0);
  signal extsi49_outs_valid : std_logic;
  signal extsi49_outs_ready : std_logic;
  signal source8_outs_valid : std_logic;
  signal source8_outs_ready : std_logic;
  signal constant43_outs : std_logic_vector(1 downto 0);
  signal constant43_outs_valid : std_logic;
  signal constant43_outs_ready : std_logic;
  signal extsi50_outs : std_logic_vector(5 downto 0);
  signal extsi50_outs_valid : std_logic;
  signal extsi50_outs_ready : std_logic;
  signal addi15_result : std_logic_vector(5 downto 0);
  signal addi15_result_valid : std_logic;
  signal addi15_result_ready : std_logic;
  signal buffer109_outs : std_logic_vector(5 downto 0);
  signal buffer109_outs_valid : std_logic;
  signal buffer109_outs_ready : std_logic;
  signal fork29_outs_0 : std_logic_vector(5 downto 0);
  signal fork29_outs_0_valid : std_logic;
  signal fork29_outs_0_ready : std_logic;
  signal fork29_outs_1 : std_logic_vector(5 downto 0);
  signal fork29_outs_1_valid : std_logic;
  signal fork29_outs_1_ready : std_logic;
  signal trunci10_outs : std_logic_vector(4 downto 0);
  signal trunci10_outs_valid : std_logic;
  signal trunci10_outs_ready : std_logic;
  signal cmpi2_result : std_logic_vector(0 downto 0);
  signal cmpi2_result_valid : std_logic;
  signal cmpi2_result_ready : std_logic;
  signal buffer114_outs : std_logic_vector(0 downto 0);
  signal buffer114_outs_valid : std_logic;
  signal buffer114_outs_ready : std_logic;
  signal fork30_outs_0 : std_logic_vector(0 downto 0);
  signal fork30_outs_0_valid : std_logic;
  signal fork30_outs_0_ready : std_logic;
  signal fork30_outs_1 : std_logic_vector(0 downto 0);
  signal fork30_outs_1_valid : std_logic;
  signal fork30_outs_1_ready : std_logic;
  signal fork30_outs_2 : std_logic_vector(0 downto 0);
  signal fork30_outs_2_valid : std_logic;
  signal fork30_outs_2_ready : std_logic;
  signal fork30_outs_3 : std_logic_vector(0 downto 0);
  signal fork30_outs_3_valid : std_logic;
  signal fork30_outs_3_ready : std_logic;
  signal fork30_outs_4 : std_logic_vector(0 downto 0);
  signal fork30_outs_4_valid : std_logic;
  signal fork30_outs_4_ready : std_logic;
  signal fork30_outs_5 : std_logic_vector(0 downto 0);
  signal fork30_outs_5_valid : std_logic;
  signal fork30_outs_5_ready : std_logic;
  signal fork30_outs_6 : std_logic_vector(0 downto 0);
  signal fork30_outs_6_valid : std_logic;
  signal fork30_outs_6_ready : std_logic;
  signal fork30_outs_7 : std_logic_vector(0 downto 0);
  signal fork30_outs_7_valid : std_logic;
  signal fork30_outs_7_ready : std_logic;
  signal cond_br17_trueOut : std_logic_vector(4 downto 0);
  signal cond_br17_trueOut_valid : std_logic;
  signal cond_br17_trueOut_ready : std_logic;
  signal cond_br17_falseOut : std_logic_vector(4 downto 0);
  signal cond_br17_falseOut_valid : std_logic;
  signal cond_br17_falseOut_ready : std_logic;
  signal cond_br18_trueOut : std_logic_vector(31 downto 0);
  signal cond_br18_trueOut_valid : std_logic;
  signal cond_br18_trueOut_ready : std_logic;
  signal cond_br18_falseOut : std_logic_vector(31 downto 0);
  signal cond_br18_falseOut_valid : std_logic;
  signal cond_br18_falseOut_ready : std_logic;
  signal cond_br19_trueOut : std_logic_vector(31 downto 0);
  signal cond_br19_trueOut_valid : std_logic;
  signal cond_br19_trueOut_ready : std_logic;
  signal cond_br19_falseOut : std_logic_vector(31 downto 0);
  signal cond_br19_falseOut_valid : std_logic;
  signal cond_br19_falseOut_ready : std_logic;
  signal cond_br20_trueOut_valid : std_logic;
  signal cond_br20_trueOut_ready : std_logic;
  signal cond_br20_falseOut_valid : std_logic;
  signal cond_br20_falseOut_ready : std_logic;
  signal cond_br21_trueOut : std_logic_vector(0 downto 0);
  signal cond_br21_trueOut_valid : std_logic;
  signal cond_br21_trueOut_ready : std_logic;
  signal cond_br21_falseOut : std_logic_vector(0 downto 0);
  signal cond_br21_falseOut_valid : std_logic;
  signal cond_br21_falseOut_ready : std_logic;
  signal extsi31_outs : std_logic_vector(4 downto 0);
  signal extsi31_outs_valid : std_logic;
  signal extsi31_outs_ready : std_logic;
  signal init14_outs : std_logic_vector(0 downto 0);
  signal init14_outs_valid : std_logic;
  signal init14_outs_ready : std_logic;
  signal fork31_outs_0 : std_logic_vector(0 downto 0);
  signal fork31_outs_0_valid : std_logic;
  signal fork31_outs_0_ready : std_logic;
  signal fork31_outs_1 : std_logic_vector(0 downto 0);
  signal fork31_outs_1_valid : std_logic;
  signal fork31_outs_1_ready : std_logic;
  signal fork31_outs_2 : std_logic_vector(0 downto 0);
  signal fork31_outs_2_valid : std_logic;
  signal fork31_outs_2_ready : std_logic;
  signal buffer215_outs_valid : std_logic;
  signal buffer215_outs_ready : std_logic;
  signal mux35_outs_valid : std_logic;
  signal mux35_outs_ready : std_logic;
  signal buffer89_outs : std_logic_vector(0 downto 0);
  signal buffer89_outs_valid : std_logic;
  signal buffer89_outs_ready : std_logic;
  signal buffer115_outs_valid : std_logic;
  signal buffer115_outs_ready : std_logic;
  signal fork32_outs_0_valid : std_logic;
  signal fork32_outs_0_ready : std_logic;
  signal fork32_outs_1_valid : std_logic;
  signal fork32_outs_1_ready : std_logic;
  signal mux36_outs_valid : std_logic;
  signal mux36_outs_ready : std_logic;
  signal buffer90_outs : std_logic_vector(0 downto 0);
  signal buffer90_outs_valid : std_logic;
  signal buffer90_outs_ready : std_logic;
  signal buffer116_outs_valid : std_logic;
  signal buffer116_outs_ready : std_logic;
  signal buffer117_outs_valid : std_logic;
  signal buffer117_outs_ready : std_logic;
  signal fork33_outs_0_valid : std_logic;
  signal fork33_outs_0_ready : std_logic;
  signal fork33_outs_1_valid : std_logic;
  signal fork33_outs_1_ready : std_logic;
  signal mux40_outs_valid : std_logic;
  signal mux40_outs_ready : std_logic;
  signal buffer91_outs : std_logic_vector(0 downto 0);
  signal buffer91_outs_valid : std_logic;
  signal buffer91_outs_ready : std_logic;
  signal mux12_outs : std_logic_vector(4 downto 0);
  signal mux12_outs_valid : std_logic;
  signal mux12_outs_ready : std_logic;
  signal mux13_outs : std_logic_vector(31 downto 0);
  signal mux13_outs_valid : std_logic;
  signal mux13_outs_ready : std_logic;
  signal control_merge5_outs_valid : std_logic;
  signal control_merge5_outs_ready : std_logic;
  signal control_merge5_index : std_logic_vector(0 downto 0);
  signal control_merge5_index_valid : std_logic;
  signal control_merge5_index_ready : std_logic;
  signal fork34_outs_0 : std_logic_vector(0 downto 0);
  signal fork34_outs_0_valid : std_logic;
  signal fork34_outs_0_ready : std_logic;
  signal fork34_outs_1 : std_logic_vector(0 downto 0);
  signal fork34_outs_1_valid : std_logic;
  signal fork34_outs_1_ready : std_logic;
  signal fork35_outs_0_valid : std_logic;
  signal fork35_outs_0_ready : std_logic;
  signal fork35_outs_1_valid : std_logic;
  signal fork35_outs_1_ready : std_logic;
  signal constant44_outs : std_logic_vector(0 downto 0);
  signal constant44_outs_valid : std_logic;
  signal constant44_outs_ready : std_logic;
  signal extsi30_outs : std_logic_vector(4 downto 0);
  signal extsi30_outs_valid : std_logic;
  signal extsi30_outs_ready : std_logic;
  signal buffer129_outs : std_logic_vector(31 downto 0);
  signal buffer129_outs_valid : std_logic;
  signal buffer129_outs_ready : std_logic;
  signal buffer130_outs : std_logic_vector(31 downto 0);
  signal buffer130_outs_valid : std_logic;
  signal buffer130_outs_ready : std_logic;
  signal buffer123_outs : std_logic_vector(4 downto 0);
  signal buffer123_outs_valid : std_logic;
  signal buffer123_outs_ready : std_logic;
  signal init20_outs : std_logic_vector(0 downto 0);
  signal init20_outs_valid : std_logic;
  signal init20_outs_ready : std_logic;
  signal fork36_outs_0 : std_logic_vector(0 downto 0);
  signal fork36_outs_0_valid : std_logic;
  signal fork36_outs_0_ready : std_logic;
  signal fork36_outs_1 : std_logic_vector(0 downto 0);
  signal fork36_outs_1_valid : std_logic;
  signal fork36_outs_1_ready : std_logic;
  signal fork36_outs_2 : std_logic_vector(0 downto 0);
  signal fork36_outs_2_valid : std_logic;
  signal fork36_outs_2_ready : std_logic;
  signal mux41_outs_valid : std_logic;
  signal mux41_outs_ready : std_logic;
  signal buffer95_outs : std_logic_vector(0 downto 0);
  signal buffer95_outs_valid : std_logic;
  signal buffer95_outs_ready : std_logic;
  signal buffer131_outs_valid : std_logic;
  signal buffer131_outs_ready : std_logic;
  signal buffer132_outs_valid : std_logic;
  signal buffer132_outs_ready : std_logic;
  signal fork37_outs_0_valid : std_logic;
  signal fork37_outs_0_ready : std_logic;
  signal fork37_outs_1_valid : std_logic;
  signal fork37_outs_1_ready : std_logic;
  signal mux42_outs_valid : std_logic;
  signal mux42_outs_ready : std_logic;
  signal buffer96_outs : std_logic_vector(0 downto 0);
  signal buffer96_outs_valid : std_logic;
  signal buffer96_outs_ready : std_logic;
  signal buffer133_outs_valid : std_logic;
  signal buffer133_outs_ready : std_logic;
  signal buffer135_outs_valid : std_logic;
  signal buffer135_outs_ready : std_logic;
  signal fork38_outs_0_valid : std_logic;
  signal fork38_outs_0_ready : std_logic;
  signal fork38_outs_1_valid : std_logic;
  signal fork38_outs_1_ready : std_logic;
  signal buffer121_outs_valid : std_logic;
  signal buffer121_outs_ready : std_logic;
  signal mux46_outs_valid : std_logic;
  signal mux46_outs_ready : std_logic;
  signal buffer97_outs : std_logic_vector(0 downto 0);
  signal buffer97_outs_valid : std_logic;
  signal buffer97_outs_ready : std_logic;
  signal unbundle2_outs_0_valid : std_logic;
  signal unbundle2_outs_0_ready : std_logic;
  signal unbundle2_outs_1 : std_logic_vector(31 downto 0);
  signal buffer98_outs : std_logic_vector(31 downto 0);
  signal buffer98_outs_valid : std_logic;
  signal buffer98_outs_ready : std_logic;
  signal mux14_outs : std_logic_vector(4 downto 0);
  signal mux14_outs_valid : std_logic;
  signal mux14_outs_ready : std_logic;
  signal buffer142_outs : std_logic_vector(4 downto 0);
  signal buffer142_outs_valid : std_logic;
  signal buffer142_outs_ready : std_logic;
  signal fork39_outs_0 : std_logic_vector(4 downto 0);
  signal fork39_outs_0_valid : std_logic;
  signal fork39_outs_0_ready : std_logic;
  signal fork39_outs_1 : std_logic_vector(4 downto 0);
  signal fork39_outs_1_valid : std_logic;
  signal fork39_outs_1_ready : std_logic;
  signal fork39_outs_2 : std_logic_vector(4 downto 0);
  signal fork39_outs_2_valid : std_logic;
  signal fork39_outs_2_ready : std_logic;
  signal extsi51_outs : std_logic_vector(6 downto 0);
  signal extsi51_outs_valid : std_logic;
  signal extsi51_outs_ready : std_logic;
  signal extsi52_outs : std_logic_vector(6 downto 0);
  signal extsi52_outs_valid : std_logic;
  signal extsi52_outs_ready : std_logic;
  signal buffer101_outs : std_logic_vector(4 downto 0);
  signal buffer101_outs_valid : std_logic;
  signal buffer101_outs_ready : std_logic;
  signal mux15_outs : std_logic_vector(31 downto 0);
  signal mux15_outs_valid : std_logic;
  signal mux15_outs_ready : std_logic;
  signal buffer145_outs : std_logic_vector(31 downto 0);
  signal buffer145_outs_valid : std_logic;
  signal buffer145_outs_ready : std_logic;
  signal fork40_outs_0 : std_logic_vector(31 downto 0);
  signal fork40_outs_0_valid : std_logic;
  signal fork40_outs_0_ready : std_logic;
  signal fork40_outs_1 : std_logic_vector(31 downto 0);
  signal fork40_outs_1_valid : std_logic;
  signal fork40_outs_1_ready : std_logic;
  signal mux16_outs : std_logic_vector(4 downto 0);
  signal mux16_outs_valid : std_logic;
  signal mux16_outs_ready : std_logic;
  signal buffer147_outs : std_logic_vector(4 downto 0);
  signal buffer147_outs_valid : std_logic;
  signal buffer147_outs_ready : std_logic;
  signal buffer161_outs : std_logic_vector(4 downto 0);
  signal buffer161_outs_valid : std_logic;
  signal buffer161_outs_ready : std_logic;
  signal fork41_outs_0 : std_logic_vector(4 downto 0);
  signal fork41_outs_0_valid : std_logic;
  signal fork41_outs_0_ready : std_logic;
  signal fork41_outs_1 : std_logic_vector(4 downto 0);
  signal fork41_outs_1_valid : std_logic;
  signal fork41_outs_1_ready : std_logic;
  signal extsi53_outs : std_logic_vector(31 downto 0);
  signal extsi53_outs_valid : std_logic;
  signal extsi53_outs_ready : std_logic;
  signal fork42_outs_0 : std_logic_vector(31 downto 0);
  signal fork42_outs_0_valid : std_logic;
  signal fork42_outs_0_ready : std_logic;
  signal fork42_outs_1 : std_logic_vector(31 downto 0);
  signal fork42_outs_1_valid : std_logic;
  signal fork42_outs_1_ready : std_logic;
  signal fork42_outs_2 : std_logic_vector(31 downto 0);
  signal fork42_outs_2_valid : std_logic;
  signal fork42_outs_2_ready : std_logic;
  signal fork42_outs_3 : std_logic_vector(31 downto 0);
  signal fork42_outs_3_valid : std_logic;
  signal fork42_outs_3_ready : std_logic;
  signal control_merge6_outs_valid : std_logic;
  signal control_merge6_outs_ready : std_logic;
  signal control_merge6_index : std_logic_vector(0 downto 0);
  signal control_merge6_index_valid : std_logic;
  signal control_merge6_index_ready : std_logic;
  signal fork43_outs_0 : std_logic_vector(0 downto 0);
  signal fork43_outs_0_valid : std_logic;
  signal fork43_outs_0_ready : std_logic;
  signal fork43_outs_1 : std_logic_vector(0 downto 0);
  signal fork43_outs_1_valid : std_logic;
  signal fork43_outs_1_ready : std_logic;
  signal fork43_outs_2 : std_logic_vector(0 downto 0);
  signal fork43_outs_2_valid : std_logic;
  signal fork43_outs_2_ready : std_logic;
  signal fork44_outs_0_valid : std_logic;
  signal fork44_outs_0_ready : std_logic;
  signal fork44_outs_1_valid : std_logic;
  signal fork44_outs_1_ready : std_logic;
  signal fork44_outs_2_valid : std_logic;
  signal fork44_outs_2_ready : std_logic;
  signal constant45_outs : std_logic_vector(1 downto 0);
  signal constant45_outs_valid : std_logic;
  signal constant45_outs_ready : std_logic;
  signal extsi17_outs : std_logic_vector(31 downto 0);
  signal extsi17_outs_valid : std_logic;
  signal extsi17_outs_ready : std_logic;
  signal constant46_outs : std_logic_vector(0 downto 0);
  signal constant46_outs_valid : std_logic;
  signal constant46_outs_ready : std_logic;
  signal source9_outs_valid : std_logic;
  signal source9_outs_ready : std_logic;
  signal constant47_outs : std_logic_vector(1 downto 0);
  signal constant47_outs_valid : std_logic;
  signal constant47_outs_ready : std_logic;
  signal extsi19_outs : std_logic_vector(31 downto 0);
  signal extsi19_outs_valid : std_logic;
  signal extsi19_outs_ready : std_logic;
  signal fork45_outs_0 : std_logic_vector(31 downto 0);
  signal fork45_outs_0_valid : std_logic;
  signal fork45_outs_0_ready : std_logic;
  signal fork45_outs_1 : std_logic_vector(31 downto 0);
  signal fork45_outs_1_valid : std_logic;
  signal fork45_outs_1_ready : std_logic;
  signal source10_outs_valid : std_logic;
  signal source10_outs_ready : std_logic;
  signal constant48_outs : std_logic_vector(2 downto 0);
  signal constant48_outs_valid : std_logic;
  signal constant48_outs_ready : std_logic;
  signal extsi20_outs : std_logic_vector(31 downto 0);
  signal extsi20_outs_valid : std_logic;
  signal extsi20_outs_ready : std_logic;
  signal fork46_outs_0 : std_logic_vector(31 downto 0);
  signal fork46_outs_0_valid : std_logic;
  signal fork46_outs_0_ready : std_logic;
  signal fork46_outs_1 : std_logic_vector(31 downto 0);
  signal fork46_outs_1_valid : std_logic;
  signal fork46_outs_1_ready : std_logic;
  signal shli10_result : std_logic_vector(31 downto 0);
  signal shli10_result_valid : std_logic;
  signal shli10_result_ready : std_logic;
  signal buffer163_outs : std_logic_vector(31 downto 0);
  signal buffer163_outs_valid : std_logic;
  signal buffer163_outs_ready : std_logic;
  signal trunci11_outs : std_logic_vector(6 downto 0);
  signal trunci11_outs_valid : std_logic;
  signal trunci11_outs_ready : std_logic;
  signal shli11_result : std_logic_vector(31 downto 0);
  signal shli11_result_valid : std_logic;
  signal shli11_result_ready : std_logic;
  signal buffer165_outs : std_logic_vector(31 downto 0);
  signal buffer165_outs_valid : std_logic;
  signal buffer165_outs_ready : std_logic;
  signal trunci12_outs : std_logic_vector(6 downto 0);
  signal trunci12_outs_valid : std_logic;
  signal trunci12_outs_ready : std_logic;
  signal addi24_result : std_logic_vector(6 downto 0);
  signal addi24_result_valid : std_logic;
  signal addi24_result_ready : std_logic;
  signal buffer168_outs : std_logic_vector(6 downto 0);
  signal buffer168_outs_valid : std_logic;
  signal buffer168_outs_ready : std_logic;
  signal addi7_result : std_logic_vector(6 downto 0);
  signal addi7_result_valid : std_logic;
  signal addi7_result_ready : std_logic;
  signal buffer2_outs_valid : std_logic;
  signal buffer2_outs_ready : std_logic;
  signal load3_addrOut : std_logic_vector(6 downto 0);
  signal load3_addrOut_valid : std_logic;
  signal load3_addrOut_ready : std_logic;
  signal load3_dataOut : std_logic_vector(31 downto 0);
  signal load3_dataOut_valid : std_logic;
  signal load3_dataOut_ready : std_logic;
  signal fork47_outs_0 : std_logic_vector(31 downto 0);
  signal fork47_outs_0_valid : std_logic;
  signal fork47_outs_0_ready : std_logic;
  signal fork47_outs_1 : std_logic_vector(31 downto 0);
  signal fork47_outs_1_valid : std_logic;
  signal fork47_outs_1_ready : std_logic;
  signal muli2_result : std_logic_vector(31 downto 0);
  signal muli2_result_valid : std_logic;
  signal muli2_result_ready : std_logic;
  signal buffer110_outs : std_logic_vector(31 downto 0);
  signal buffer110_outs_valid : std_logic;
  signal buffer110_outs_ready : std_logic;
  signal shli12_result : std_logic_vector(31 downto 0);
  signal shli12_result_valid : std_logic;
  signal shli12_result_ready : std_logic;
  signal buffer111_outs : std_logic_vector(31 downto 0);
  signal buffer111_outs_valid : std_logic;
  signal buffer111_outs_ready : std_logic;
  signal buffer112_outs : std_logic_vector(31 downto 0);
  signal buffer112_outs_valid : std_logic;
  signal buffer112_outs_ready : std_logic;
  signal buffer171_outs : std_logic_vector(31 downto 0);
  signal buffer171_outs_valid : std_logic;
  signal buffer171_outs_ready : std_logic;
  signal trunci13_outs : std_logic_vector(6 downto 0);
  signal trunci13_outs_valid : std_logic;
  signal trunci13_outs_ready : std_logic;
  signal shli13_result : std_logic_vector(31 downto 0);
  signal shli13_result_valid : std_logic;
  signal shli13_result_ready : std_logic;
  signal buffer113_outs : std_logic_vector(31 downto 0);
  signal buffer113_outs_valid : std_logic;
  signal buffer113_outs_ready : std_logic;
  signal buffer172_outs : std_logic_vector(31 downto 0);
  signal buffer172_outs_valid : std_logic;
  signal buffer172_outs_ready : std_logic;
  signal trunci14_outs : std_logic_vector(6 downto 0);
  signal trunci14_outs_valid : std_logic;
  signal trunci14_outs_ready : std_logic;
  signal addi25_result : std_logic_vector(6 downto 0);
  signal addi25_result_valid : std_logic;
  signal addi25_result_ready : std_logic;
  signal buffer173_outs : std_logic_vector(6 downto 0);
  signal buffer173_outs_valid : std_logic;
  signal buffer173_outs_ready : std_logic;
  signal addi8_result : std_logic_vector(6 downto 0);
  signal addi8_result_valid : std_logic;
  signal addi8_result_ready : std_logic;
  signal buffer3_outs_valid : std_logic;
  signal buffer3_outs_ready : std_logic;
  signal buffer175_outs : std_logic_vector(6 downto 0);
  signal buffer175_outs_valid : std_logic;
  signal buffer175_outs_ready : std_logic;
  signal store2_addrOut : std_logic_vector(6 downto 0);
  signal store2_addrOut_valid : std_logic;
  signal store2_addrOut_ready : std_logic;
  signal store2_dataToMem : std_logic_vector(31 downto 0);
  signal store2_dataToMem_valid : std_logic;
  signal store2_dataToMem_ready : std_logic;
  signal store2_doneOut_valid : std_logic;
  signal store2_doneOut_ready : std_logic;
  signal extsi29_outs : std_logic_vector(4 downto 0);
  signal extsi29_outs_valid : std_logic;
  signal extsi29_outs_ready : std_logic;
  signal cond_br89_trueOut_valid : std_logic;
  signal cond_br89_trueOut_ready : std_logic;
  signal cond_br89_falseOut_valid : std_logic;
  signal cond_br89_falseOut_ready : std_logic;
  signal buffer118_outs : std_logic_vector(0 downto 0);
  signal buffer118_outs_valid : std_logic;
  signal buffer118_outs_ready : std_logic;
  signal cond_br90_trueOut_valid : std_logic;
  signal cond_br90_trueOut_ready : std_logic;
  signal cond_br90_falseOut_valid : std_logic;
  signal cond_br90_falseOut_ready : std_logic;
  signal buffer119_outs : std_logic_vector(0 downto 0);
  signal buffer119_outs_valid : std_logic;
  signal buffer119_outs_ready : std_logic;
  signal cond_br91_trueOut_valid : std_logic;
  signal cond_br91_trueOut_ready : std_logic;
  signal cond_br91_falseOut_valid : std_logic;
  signal cond_br91_falseOut_ready : std_logic;
  signal buffer120_outs : std_logic_vector(0 downto 0);
  signal buffer120_outs_valid : std_logic;
  signal buffer120_outs_ready : std_logic;
  signal cond_br92_trueOut_valid : std_logic;
  signal cond_br92_trueOut_ready : std_logic;
  signal cond_br92_falseOut_valid : std_logic;
  signal cond_br92_falseOut_ready : std_logic;
  signal buffer209_outs_valid : std_logic;
  signal buffer209_outs_ready : std_logic;
  signal cond_br93_trueOut_valid : std_logic;
  signal cond_br93_trueOut_ready : std_logic;
  signal cond_br93_falseOut_valid : std_logic;
  signal cond_br93_falseOut_ready : std_logic;
  signal buffer122_outs : std_logic_vector(0 downto 0);
  signal buffer122_outs_valid : std_logic;
  signal buffer122_outs_ready : std_logic;
  signal init26_outs : std_logic_vector(0 downto 0);
  signal init26_outs_valid : std_logic;
  signal init26_outs_ready : std_logic;
  signal fork48_outs_0 : std_logic_vector(0 downto 0);
  signal fork48_outs_0_valid : std_logic;
  signal fork48_outs_0_ready : std_logic;
  signal fork48_outs_1 : std_logic_vector(0 downto 0);
  signal fork48_outs_1_valid : std_logic;
  signal fork48_outs_1_ready : std_logic;
  signal fork48_outs_2 : std_logic_vector(0 downto 0);
  signal fork48_outs_2_valid : std_logic;
  signal fork48_outs_2_ready : std_logic;
  signal fork48_outs_3 : std_logic_vector(0 downto 0);
  signal fork48_outs_3_valid : std_logic;
  signal fork48_outs_3_ready : std_logic;
  signal fork48_outs_4 : std_logic_vector(0 downto 0);
  signal fork48_outs_4_valid : std_logic;
  signal fork48_outs_4_ready : std_logic;
  signal mux47_outs_valid : std_logic;
  signal mux47_outs_ready : std_logic;
  signal buffer124_outs : std_logic_vector(0 downto 0);
  signal buffer124_outs_valid : std_logic;
  signal buffer124_outs_ready : std_logic;
  signal buffer178_outs_valid : std_logic;
  signal buffer178_outs_ready : std_logic;
  signal buffer179_outs_valid : std_logic;
  signal buffer179_outs_ready : std_logic;
  signal fork49_outs_0_valid : std_logic;
  signal fork49_outs_0_ready : std_logic;
  signal fork49_outs_1_valid : std_logic;
  signal fork49_outs_1_ready : std_logic;
  signal fork49_outs_2_valid : std_logic;
  signal fork49_outs_2_ready : std_logic;
  signal mux48_outs_valid : std_logic;
  signal mux48_outs_ready : std_logic;
  signal buffer125_outs : std_logic_vector(0 downto 0);
  signal buffer125_outs_valid : std_logic;
  signal buffer125_outs_ready : std_logic;
  signal buffer180_outs_valid : std_logic;
  signal buffer180_outs_ready : std_logic;
  signal buffer181_outs_valid : std_logic;
  signal buffer181_outs_ready : std_logic;
  signal fork50_outs_0_valid : std_logic;
  signal fork50_outs_0_ready : std_logic;
  signal fork50_outs_1_valid : std_logic;
  signal fork50_outs_1_ready : std_logic;
  signal mux49_outs_valid : std_logic;
  signal mux49_outs_ready : std_logic;
  signal buffer126_outs : std_logic_vector(0 downto 0);
  signal buffer126_outs_valid : std_logic;
  signal buffer126_outs_ready : std_logic;
  signal buffer182_outs_valid : std_logic;
  signal buffer182_outs_ready : std_logic;
  signal buffer183_outs_valid : std_logic;
  signal buffer183_outs_ready : std_logic;
  signal fork51_outs_0_valid : std_logic;
  signal fork51_outs_0_ready : std_logic;
  signal fork51_outs_1_valid : std_logic;
  signal fork51_outs_1_ready : std_logic;
  signal mux51_outs_valid : std_logic;
  signal mux51_outs_ready : std_logic;
  signal buffer127_outs : std_logic_vector(0 downto 0);
  signal buffer127_outs_valid : std_logic;
  signal buffer127_outs_ready : std_logic;
  signal buffer185_outs_valid : std_logic;
  signal buffer185_outs_ready : std_logic;
  signal buffer186_outs_valid : std_logic;
  signal buffer186_outs_ready : std_logic;
  signal fork52_outs_0_valid : std_logic;
  signal fork52_outs_0_ready : std_logic;
  signal fork52_outs_1_valid : std_logic;
  signal fork52_outs_1_ready : std_logic;
  signal buffer136_outs_valid : std_logic;
  signal buffer136_outs_ready : std_logic;
  signal buffer140_outs_valid : std_logic;
  signal buffer140_outs_ready : std_logic;
  signal mux52_outs_valid : std_logic;
  signal mux52_outs_ready : std_logic;
  signal buffer128_outs : std_logic_vector(0 downto 0);
  signal buffer128_outs_valid : std_logic;
  signal buffer128_outs_ready : std_logic;
  signal mux17_outs : std_logic_vector(4 downto 0);
  signal mux17_outs_valid : std_logic;
  signal mux17_outs_ready : std_logic;
  signal buffer188_outs : std_logic_vector(4 downto 0);
  signal buffer188_outs_valid : std_logic;
  signal buffer188_outs_ready : std_logic;
  signal buffer189_outs : std_logic_vector(4 downto 0);
  signal buffer189_outs_valid : std_logic;
  signal buffer189_outs_ready : std_logic;
  signal fork53_outs_0 : std_logic_vector(4 downto 0);
  signal fork53_outs_0_valid : std_logic;
  signal fork53_outs_0_ready : std_logic;
  signal fork53_outs_1 : std_logic_vector(4 downto 0);
  signal fork53_outs_1_valid : std_logic;
  signal fork53_outs_1_ready : std_logic;
  signal extsi54_outs : std_logic_vector(5 downto 0);
  signal extsi54_outs_valid : std_logic;
  signal extsi54_outs_ready : std_logic;
  signal extsi55_outs : std_logic_vector(31 downto 0);
  signal extsi55_outs_valid : std_logic;
  signal extsi55_outs_ready : std_logic;
  signal fork54_outs_0 : std_logic_vector(31 downto 0);
  signal fork54_outs_0_valid : std_logic;
  signal fork54_outs_0_ready : std_logic;
  signal fork54_outs_1 : std_logic_vector(31 downto 0);
  signal fork54_outs_1_valid : std_logic;
  signal fork54_outs_1_ready : std_logic;
  signal fork54_outs_2 : std_logic_vector(31 downto 0);
  signal fork54_outs_2_valid : std_logic;
  signal fork54_outs_2_ready : std_logic;
  signal mux18_outs : std_logic_vector(31 downto 0);
  signal mux18_outs_valid : std_logic;
  signal mux18_outs_ready : std_logic;
  signal mux19_outs : std_logic_vector(4 downto 0);
  signal mux19_outs_valid : std_logic;
  signal mux19_outs_ready : std_logic;
  signal buffer192_outs : std_logic_vector(4 downto 0);
  signal buffer192_outs_valid : std_logic;
  signal buffer192_outs_ready : std_logic;
  signal buffer193_outs : std_logic_vector(4 downto 0);
  signal buffer193_outs_valid : std_logic;
  signal buffer193_outs_ready : std_logic;
  signal fork55_outs_0 : std_logic_vector(4 downto 0);
  signal fork55_outs_0_valid : std_logic;
  signal fork55_outs_0_ready : std_logic;
  signal fork55_outs_1 : std_logic_vector(4 downto 0);
  signal fork55_outs_1_valid : std_logic;
  signal fork55_outs_1_ready : std_logic;
  signal extsi56_outs : std_logic_vector(31 downto 0);
  signal extsi56_outs_valid : std_logic;
  signal extsi56_outs_ready : std_logic;
  signal buffer134_outs : std_logic_vector(4 downto 0);
  signal buffer134_outs_valid : std_logic;
  signal buffer134_outs_ready : std_logic;
  signal fork56_outs_0 : std_logic_vector(31 downto 0);
  signal fork56_outs_0_valid : std_logic;
  signal fork56_outs_0_ready : std_logic;
  signal fork56_outs_1 : std_logic_vector(31 downto 0);
  signal fork56_outs_1_valid : std_logic;
  signal fork56_outs_1_ready : std_logic;
  signal fork56_outs_2 : std_logic_vector(31 downto 0);
  signal fork56_outs_2_valid : std_logic;
  signal fork56_outs_2_ready : std_logic;
  signal fork56_outs_3 : std_logic_vector(31 downto 0);
  signal fork56_outs_3_valid : std_logic;
  signal fork56_outs_3_ready : std_logic;
  signal fork56_outs_4 : std_logic_vector(31 downto 0);
  signal fork56_outs_4_valid : std_logic;
  signal fork56_outs_4_ready : std_logic;
  signal fork56_outs_5 : std_logic_vector(31 downto 0);
  signal fork56_outs_5_valid : std_logic;
  signal fork56_outs_5_ready : std_logic;
  signal mux20_outs : std_logic_vector(4 downto 0);
  signal mux20_outs_valid : std_logic;
  signal mux20_outs_ready : std_logic;
  signal buffer194_outs : std_logic_vector(4 downto 0);
  signal buffer194_outs_valid : std_logic;
  signal buffer194_outs_ready : std_logic;
  signal buffer195_outs : std_logic_vector(4 downto 0);
  signal buffer195_outs_valid : std_logic;
  signal buffer195_outs_ready : std_logic;
  signal fork57_outs_0 : std_logic_vector(4 downto 0);
  signal fork57_outs_0_valid : std_logic;
  signal fork57_outs_0_ready : std_logic;
  signal fork57_outs_1 : std_logic_vector(4 downto 0);
  signal fork57_outs_1_valid : std_logic;
  signal fork57_outs_1_ready : std_logic;
  signal fork57_outs_2 : std_logic_vector(4 downto 0);
  signal fork57_outs_2_valid : std_logic;
  signal fork57_outs_2_ready : std_logic;
  signal extsi57_outs : std_logic_vector(6 downto 0);
  signal extsi57_outs_valid : std_logic;
  signal extsi57_outs_ready : std_logic;
  signal extsi58_outs : std_logic_vector(31 downto 0);
  signal extsi58_outs_valid : std_logic;
  signal extsi58_outs_ready : std_logic;
  signal buffer137_outs : std_logic_vector(4 downto 0);
  signal buffer137_outs_valid : std_logic;
  signal buffer137_outs_ready : std_logic;
  signal fork58_outs_0 : std_logic_vector(31 downto 0);
  signal fork58_outs_0_valid : std_logic;
  signal fork58_outs_0_ready : std_logic;
  signal fork58_outs_1 : std_logic_vector(31 downto 0);
  signal fork58_outs_1_valid : std_logic;
  signal fork58_outs_1_ready : std_logic;
  signal control_merge7_outs_valid : std_logic;
  signal control_merge7_outs_ready : std_logic;
  signal control_merge7_index : std_logic_vector(0 downto 0);
  signal control_merge7_index_valid : std_logic;
  signal control_merge7_index_ready : std_logic;
  signal fork59_outs_0 : std_logic_vector(0 downto 0);
  signal fork59_outs_0_valid : std_logic;
  signal fork59_outs_0_ready : std_logic;
  signal fork59_outs_1 : std_logic_vector(0 downto 0);
  signal fork59_outs_1_valid : std_logic;
  signal fork59_outs_1_ready : std_logic;
  signal fork59_outs_2 : std_logic_vector(0 downto 0);
  signal fork59_outs_2_valid : std_logic;
  signal fork59_outs_2_ready : std_logic;
  signal fork59_outs_3 : std_logic_vector(0 downto 0);
  signal fork59_outs_3_valid : std_logic;
  signal fork59_outs_3_ready : std_logic;
  signal buffer196_outs_valid : std_logic;
  signal buffer196_outs_ready : std_logic;
  signal fork60_outs_0_valid : std_logic;
  signal fork60_outs_0_ready : std_logic;
  signal fork60_outs_1_valid : std_logic;
  signal fork60_outs_1_ready : std_logic;
  signal constant49_outs : std_logic_vector(1 downto 0);
  signal constant49_outs_valid : std_logic;
  signal constant49_outs_ready : std_logic;
  signal extsi21_outs : std_logic_vector(31 downto 0);
  signal extsi21_outs_valid : std_logic;
  signal extsi21_outs_ready : std_logic;
  signal source11_outs_valid : std_logic;
  signal source11_outs_ready : std_logic;
  signal constant50_outs : std_logic_vector(4 downto 0);
  signal constant50_outs_valid : std_logic;
  signal constant50_outs_ready : std_logic;
  signal extsi59_outs : std_logic_vector(5 downto 0);
  signal extsi59_outs_valid : std_logic;
  signal extsi59_outs_ready : std_logic;
  signal source12_outs_valid : std_logic;
  signal source12_outs_ready : std_logic;
  signal constant51_outs : std_logic_vector(1 downto 0);
  signal constant51_outs_valid : std_logic;
  signal constant51_outs_ready : std_logic;
  signal fork61_outs_0 : std_logic_vector(1 downto 0);
  signal fork61_outs_0_valid : std_logic;
  signal fork61_outs_0_ready : std_logic;
  signal fork61_outs_1 : std_logic_vector(1 downto 0);
  signal fork61_outs_1_valid : std_logic;
  signal fork61_outs_1_ready : std_logic;
  signal extsi60_outs : std_logic_vector(5 downto 0);
  signal extsi60_outs_valid : std_logic;
  signal extsi60_outs_ready : std_logic;
  signal buffer138_outs : std_logic_vector(1 downto 0);
  signal buffer138_outs_valid : std_logic;
  signal buffer138_outs_ready : std_logic;
  signal extsi23_outs : std_logic_vector(31 downto 0);
  signal extsi23_outs_valid : std_logic;
  signal extsi23_outs_ready : std_logic;
  signal buffer139_outs : std_logic_vector(1 downto 0);
  signal buffer139_outs_valid : std_logic;
  signal buffer139_outs_ready : std_logic;
  signal fork62_outs_0 : std_logic_vector(31 downto 0);
  signal fork62_outs_0_valid : std_logic;
  signal fork62_outs_0_ready : std_logic;
  signal fork62_outs_1 : std_logic_vector(31 downto 0);
  signal fork62_outs_1_valid : std_logic;
  signal fork62_outs_1_ready : std_logic;
  signal fork62_outs_2 : std_logic_vector(31 downto 0);
  signal fork62_outs_2_valid : std_logic;
  signal fork62_outs_2_ready : std_logic;
  signal fork62_outs_3 : std_logic_vector(31 downto 0);
  signal fork62_outs_3_valid : std_logic;
  signal fork62_outs_3_ready : std_logic;
  signal source13_outs_valid : std_logic;
  signal source13_outs_ready : std_logic;
  signal constant52_outs : std_logic_vector(2 downto 0);
  signal constant52_outs_valid : std_logic;
  signal constant52_outs_ready : std_logic;
  signal extsi24_outs : std_logic_vector(31 downto 0);
  signal extsi24_outs_valid : std_logic;
  signal extsi24_outs_ready : std_logic;
  signal fork63_outs_0 : std_logic_vector(31 downto 0);
  signal fork63_outs_0_valid : std_logic;
  signal fork63_outs_0_ready : std_logic;
  signal fork63_outs_1 : std_logic_vector(31 downto 0);
  signal fork63_outs_1_valid : std_logic;
  signal fork63_outs_1_ready : std_logic;
  signal fork63_outs_2 : std_logic_vector(31 downto 0);
  signal fork63_outs_2_valid : std_logic;
  signal fork63_outs_2_ready : std_logic;
  signal fork63_outs_3 : std_logic_vector(31 downto 0);
  signal fork63_outs_3_valid : std_logic;
  signal fork63_outs_3_ready : std_logic;
  signal shli14_result : std_logic_vector(31 downto 0);
  signal shli14_result_valid : std_logic;
  signal shli14_result_ready : std_logic;
  signal buffer141_outs : std_logic_vector(31 downto 0);
  signal buffer141_outs_valid : std_logic;
  signal buffer141_outs_ready : std_logic;
  signal shli15_result : std_logic_vector(31 downto 0);
  signal shli15_result_valid : std_logic;
  signal shli15_result_ready : std_logic;
  signal buffer143_outs : std_logic_vector(31 downto 0);
  signal buffer143_outs_valid : std_logic;
  signal buffer143_outs_ready : std_logic;
  signal buffer197_outs : std_logic_vector(31 downto 0);
  signal buffer197_outs_valid : std_logic;
  signal buffer197_outs_ready : std_logic;
  signal buffer198_outs : std_logic_vector(31 downto 0);
  signal buffer198_outs_valid : std_logic;
  signal buffer198_outs_ready : std_logic;
  signal addi26_result : std_logic_vector(31 downto 0);
  signal addi26_result_valid : std_logic;
  signal addi26_result_ready : std_logic;
  signal buffer199_outs : std_logic_vector(31 downto 0);
  signal buffer199_outs_valid : std_logic;
  signal buffer199_outs_ready : std_logic;
  signal addi9_result : std_logic_vector(31 downto 0);
  signal addi9_result_valid : std_logic;
  signal addi9_result_ready : std_logic;
  signal buffer144_outs : std_logic_vector(31 downto 0);
  signal buffer144_outs_valid : std_logic;
  signal buffer144_outs_ready : std_logic;
  signal gate2_outs : std_logic_vector(31 downto 0);
  signal gate2_outs_valid : std_logic;
  signal gate2_outs_ready : std_logic;
  signal trunci15_outs : std_logic_vector(6 downto 0);
  signal trunci15_outs_valid : std_logic;
  signal trunci15_outs_ready : std_logic;
  signal load4_addrOut : std_logic_vector(6 downto 0);
  signal load4_addrOut_valid : std_logic;
  signal load4_addrOut_ready : std_logic;
  signal load4_dataOut : std_logic_vector(31 downto 0);
  signal load4_dataOut_valid : std_logic;
  signal load4_dataOut_ready : std_logic;
  signal shli16_result : std_logic_vector(31 downto 0);
  signal shli16_result_valid : std_logic;
  signal shli16_result_ready : std_logic;
  signal buffer146_outs : std_logic_vector(31 downto 0);
  signal buffer146_outs_valid : std_logic;
  signal buffer146_outs_ready : std_logic;
  signal buffer200_outs : std_logic_vector(31 downto 0);
  signal buffer200_outs_valid : std_logic;
  signal buffer200_outs_ready : std_logic;
  signal trunci16_outs : std_logic_vector(6 downto 0);
  signal trunci16_outs_valid : std_logic;
  signal trunci16_outs_ready : std_logic;
  signal shli17_result : std_logic_vector(31 downto 0);
  signal shli17_result_valid : std_logic;
  signal shli17_result_ready : std_logic;
  signal buffer148_outs : std_logic_vector(31 downto 0);
  signal buffer148_outs_valid : std_logic;
  signal buffer148_outs_ready : std_logic;
  signal buffer201_outs : std_logic_vector(31 downto 0);
  signal buffer201_outs_valid : std_logic;
  signal buffer201_outs_ready : std_logic;
  signal trunci17_outs : std_logic_vector(6 downto 0);
  signal trunci17_outs_valid : std_logic;
  signal trunci17_outs_ready : std_logic;
  signal addi27_result : std_logic_vector(6 downto 0);
  signal addi27_result_valid : std_logic;
  signal addi27_result_ready : std_logic;
  signal buffer202_outs : std_logic_vector(6 downto 0);
  signal buffer202_outs_valid : std_logic;
  signal buffer202_outs_ready : std_logic;
  signal addi10_result : std_logic_vector(6 downto 0);
  signal addi10_result_valid : std_logic;
  signal addi10_result_ready : std_logic;
  signal load5_addrOut : std_logic_vector(6 downto 0);
  signal load5_addrOut_valid : std_logic;
  signal load5_addrOut_ready : std_logic;
  signal load5_dataOut : std_logic_vector(31 downto 0);
  signal load5_dataOut_valid : std_logic;
  signal load5_dataOut_ready : std_logic;
  signal muli3_result : std_logic_vector(31 downto 0);
  signal muli3_result_valid : std_logic;
  signal muli3_result_ready : std_logic;
  signal shli18_result : std_logic_vector(31 downto 0);
  signal shli18_result_valid : std_logic;
  signal shli18_result_ready : std_logic;
  signal buffer149_outs : std_logic_vector(31 downto 0);
  signal buffer149_outs_valid : std_logic;
  signal buffer149_outs_ready : std_logic;
  signal buffer150_outs : std_logic_vector(31 downto 0);
  signal buffer150_outs_valid : std_logic;
  signal buffer150_outs_ready : std_logic;
  signal shli19_result : std_logic_vector(31 downto 0);
  signal shli19_result_valid : std_logic;
  signal shli19_result_ready : std_logic;
  signal buffer151_outs : std_logic_vector(31 downto 0);
  signal buffer151_outs_valid : std_logic;
  signal buffer151_outs_ready : std_logic;
  signal buffer152_outs : std_logic_vector(31 downto 0);
  signal buffer152_outs_valid : std_logic;
  signal buffer152_outs_ready : std_logic;
  signal buffer203_outs : std_logic_vector(31 downto 0);
  signal buffer203_outs_valid : std_logic;
  signal buffer203_outs_ready : std_logic;
  signal buffer204_outs : std_logic_vector(31 downto 0);
  signal buffer204_outs_valid : std_logic;
  signal buffer204_outs_ready : std_logic;
  signal addi28_result : std_logic_vector(31 downto 0);
  signal addi28_result_valid : std_logic;
  signal addi28_result_ready : std_logic;
  signal buffer205_outs : std_logic_vector(31 downto 0);
  signal buffer205_outs_valid : std_logic;
  signal buffer205_outs_ready : std_logic;
  signal addi11_result : std_logic_vector(31 downto 0);
  signal addi11_result_valid : std_logic;
  signal addi11_result_ready : std_logic;
  signal buffer153_outs : std_logic_vector(31 downto 0);
  signal buffer153_outs_valid : std_logic;
  signal buffer153_outs_ready : std_logic;
  signal buffer187_outs_valid : std_logic;
  signal buffer187_outs_ready : std_logic;
  signal gate3_outs : std_logic_vector(31 downto 0);
  signal gate3_outs_valid : std_logic;
  signal gate3_outs_ready : std_logic;
  signal trunci18_outs : std_logic_vector(6 downto 0);
  signal trunci18_outs_valid : std_logic;
  signal trunci18_outs_ready : std_logic;
  signal load6_addrOut : std_logic_vector(6 downto 0);
  signal load6_addrOut_valid : std_logic;
  signal load6_addrOut_ready : std_logic;
  signal load6_dataOut : std_logic_vector(31 downto 0);
  signal load6_dataOut_valid : std_logic;
  signal load6_dataOut_ready : std_logic;
  signal addi1_result : std_logic_vector(31 downto 0);
  signal addi1_result_valid : std_logic;
  signal addi1_result_ready : std_logic;
  signal shli20_result : std_logic_vector(31 downto 0);
  signal shli20_result_valid : std_logic;
  signal shli20_result_ready : std_logic;
  signal buffer154_outs : std_logic_vector(31 downto 0);
  signal buffer154_outs_valid : std_logic;
  signal buffer154_outs_ready : std_logic;
  signal buffer155_outs : std_logic_vector(31 downto 0);
  signal buffer155_outs_valid : std_logic;
  signal buffer155_outs_ready : std_logic;
  signal shli21_result : std_logic_vector(31 downto 0);
  signal shli21_result_valid : std_logic;
  signal shli21_result_ready : std_logic;
  signal buffer156_outs : std_logic_vector(31 downto 0);
  signal buffer156_outs_valid : std_logic;
  signal buffer156_outs_ready : std_logic;
  signal buffer157_outs : std_logic_vector(31 downto 0);
  signal buffer157_outs_valid : std_logic;
  signal buffer157_outs_ready : std_logic;
  signal buffer206_outs : std_logic_vector(31 downto 0);
  signal buffer206_outs_valid : std_logic;
  signal buffer206_outs_ready : std_logic;
  signal buffer207_outs : std_logic_vector(31 downto 0);
  signal buffer207_outs_valid : std_logic;
  signal buffer207_outs_ready : std_logic;
  signal addi29_result : std_logic_vector(31 downto 0);
  signal addi29_result_valid : std_logic;
  signal addi29_result_ready : std_logic;
  signal buffer208_outs : std_logic_vector(31 downto 0);
  signal buffer208_outs_valid : std_logic;
  signal buffer208_outs_ready : std_logic;
  signal addi12_result : std_logic_vector(31 downto 0);
  signal addi12_result_valid : std_logic;
  signal addi12_result_ready : std_logic;
  signal buffer158_outs : std_logic_vector(31 downto 0);
  signal buffer158_outs_valid : std_logic;
  signal buffer158_outs_ready : std_logic;
  signal buffer4_outs_valid : std_logic;
  signal buffer4_outs_ready : std_logic;
  signal gate4_outs : std_logic_vector(31 downto 0);
  signal gate4_outs_valid : std_logic;
  signal gate4_outs_ready : std_logic;
  signal trunci19_outs : std_logic_vector(6 downto 0);
  signal trunci19_outs_valid : std_logic;
  signal trunci19_outs_ready : std_logic;
  signal store3_addrOut : std_logic_vector(6 downto 0);
  signal store3_addrOut_valid : std_logic;
  signal store3_addrOut_ready : std_logic;
  signal store3_dataToMem : std_logic_vector(31 downto 0);
  signal store3_dataToMem_valid : std_logic;
  signal store3_dataToMem_ready : std_logic;
  signal store3_doneOut_valid : std_logic;
  signal store3_doneOut_ready : std_logic;
  signal addi16_result : std_logic_vector(5 downto 0);
  signal addi16_result_valid : std_logic;
  signal addi16_result_ready : std_logic;
  signal fork64_outs_0 : std_logic_vector(5 downto 0);
  signal fork64_outs_0_valid : std_logic;
  signal fork64_outs_0_ready : std_logic;
  signal fork64_outs_1 : std_logic_vector(5 downto 0);
  signal fork64_outs_1_valid : std_logic;
  signal fork64_outs_1_ready : std_logic;
  signal trunci20_outs : std_logic_vector(4 downto 0);
  signal trunci20_outs_valid : std_logic;
  signal trunci20_outs_ready : std_logic;
  signal buffer159_outs : std_logic_vector(5 downto 0);
  signal buffer159_outs_valid : std_logic;
  signal buffer159_outs_ready : std_logic;
  signal cmpi3_result : std_logic_vector(0 downto 0);
  signal cmpi3_result_valid : std_logic;
  signal cmpi3_result_ready : std_logic;
  signal buffer210_outs : std_logic_vector(5 downto 0);
  signal buffer210_outs_valid : std_logic;
  signal buffer210_outs_ready : std_logic;
  signal buffer160_outs : std_logic_vector(5 downto 0);
  signal buffer160_outs_valid : std_logic;
  signal buffer160_outs_ready : std_logic;
  signal buffer211_outs : std_logic_vector(0 downto 0);
  signal buffer211_outs_valid : std_logic;
  signal buffer211_outs_ready : std_logic;
  signal fork65_outs_0 : std_logic_vector(0 downto 0);
  signal fork65_outs_0_valid : std_logic;
  signal fork65_outs_0_ready : std_logic;
  signal fork65_outs_1 : std_logic_vector(0 downto 0);
  signal fork65_outs_1_valid : std_logic;
  signal fork65_outs_1_ready : std_logic;
  signal fork65_outs_2 : std_logic_vector(0 downto 0);
  signal fork65_outs_2_valid : std_logic;
  signal fork65_outs_2_ready : std_logic;
  signal fork65_outs_3 : std_logic_vector(0 downto 0);
  signal fork65_outs_3_valid : std_logic;
  signal fork65_outs_3_ready : std_logic;
  signal fork65_outs_4 : std_logic_vector(0 downto 0);
  signal fork65_outs_4_valid : std_logic;
  signal fork65_outs_4_ready : std_logic;
  signal fork65_outs_5 : std_logic_vector(0 downto 0);
  signal fork65_outs_5_valid : std_logic;
  signal fork65_outs_5_ready : std_logic;
  signal fork65_outs_6 : std_logic_vector(0 downto 0);
  signal fork65_outs_6_valid : std_logic;
  signal fork65_outs_6_ready : std_logic;
  signal fork65_outs_7 : std_logic_vector(0 downto 0);
  signal fork65_outs_7_valid : std_logic;
  signal fork65_outs_7_ready : std_logic;
  signal fork65_outs_8 : std_logic_vector(0 downto 0);
  signal fork65_outs_8_valid : std_logic;
  signal fork65_outs_8_ready : std_logic;
  signal fork65_outs_9 : std_logic_vector(0 downto 0);
  signal fork65_outs_9_valid : std_logic;
  signal fork65_outs_9_ready : std_logic;
  signal fork65_outs_10 : std_logic_vector(0 downto 0);
  signal fork65_outs_10_valid : std_logic;
  signal fork65_outs_10_ready : std_logic;
  signal cond_br22_trueOut : std_logic_vector(4 downto 0);
  signal cond_br22_trueOut_valid : std_logic;
  signal cond_br22_trueOut_ready : std_logic;
  signal cond_br22_falseOut : std_logic_vector(4 downto 0);
  signal cond_br22_falseOut_valid : std_logic;
  signal cond_br22_falseOut_ready : std_logic;
  signal buffer190_outs : std_logic_vector(31 downto 0);
  signal buffer190_outs_valid : std_logic;
  signal buffer190_outs_ready : std_logic;
  signal buffer191_outs : std_logic_vector(31 downto 0);
  signal buffer191_outs_valid : std_logic;
  signal buffer191_outs_ready : std_logic;
  signal cond_br23_trueOut : std_logic_vector(31 downto 0);
  signal cond_br23_trueOut_valid : std_logic;
  signal cond_br23_trueOut_ready : std_logic;
  signal cond_br23_falseOut : std_logic_vector(31 downto 0);
  signal cond_br23_falseOut_valid : std_logic;
  signal cond_br23_falseOut_ready : std_logic;
  signal buffer162_outs : std_logic_vector(0 downto 0);
  signal buffer162_outs_valid : std_logic;
  signal buffer162_outs_ready : std_logic;
  signal cond_br24_trueOut : std_logic_vector(4 downto 0);
  signal cond_br24_trueOut_valid : std_logic;
  signal cond_br24_trueOut_ready : std_logic;
  signal cond_br24_falseOut : std_logic_vector(4 downto 0);
  signal cond_br24_falseOut_valid : std_logic;
  signal cond_br24_falseOut_ready : std_logic;
  signal buffer164_outs : std_logic_vector(4 downto 0);
  signal buffer164_outs_valid : std_logic;
  signal buffer164_outs_ready : std_logic;
  signal cond_br25_trueOut : std_logic_vector(4 downto 0);
  signal cond_br25_trueOut_valid : std_logic;
  signal cond_br25_trueOut_ready : std_logic;
  signal cond_br25_falseOut : std_logic_vector(4 downto 0);
  signal cond_br25_falseOut_valid : std_logic;
  signal cond_br25_falseOut_ready : std_logic;
  signal buffer166_outs : std_logic_vector(4 downto 0);
  signal buffer166_outs_valid : std_logic;
  signal buffer166_outs_ready : std_logic;
  signal cond_br26_trueOut_valid : std_logic;
  signal cond_br26_trueOut_ready : std_logic;
  signal cond_br26_falseOut_valid : std_logic;
  signal cond_br26_falseOut_ready : std_logic;
  signal buffer167_outs : std_logic_vector(0 downto 0);
  signal buffer167_outs_valid : std_logic;
  signal buffer167_outs_ready : std_logic;
  signal cond_br94_trueOut_valid : std_logic;
  signal cond_br94_trueOut_ready : std_logic;
  signal cond_br94_falseOut_valid : std_logic;
  signal cond_br94_falseOut_ready : std_logic;
  signal cond_br95_trueOut_valid : std_logic;
  signal cond_br95_trueOut_ready : std_logic;
  signal cond_br95_falseOut_valid : std_logic;
  signal cond_br95_falseOut_ready : std_logic;
  signal buffer169_outs : std_logic_vector(0 downto 0);
  signal buffer169_outs_valid : std_logic;
  signal buffer169_outs_ready : std_logic;
  signal cond_br96_trueOut_valid : std_logic;
  signal cond_br96_trueOut_ready : std_logic;
  signal cond_br96_falseOut_valid : std_logic;
  signal cond_br96_falseOut_ready : std_logic;
  signal buffer170_outs : std_logic_vector(0 downto 0);
  signal buffer170_outs_valid : std_logic;
  signal buffer170_outs_ready : std_logic;
  signal extsi61_outs : std_logic_vector(5 downto 0);
  signal extsi61_outs_valid : std_logic;
  signal extsi61_outs_ready : std_logic;
  signal source14_outs_valid : std_logic;
  signal source14_outs_ready : std_logic;
  signal constant53_outs : std_logic_vector(4 downto 0);
  signal constant53_outs_valid : std_logic;
  signal constant53_outs_ready : std_logic;
  signal extsi62_outs : std_logic_vector(5 downto 0);
  signal extsi62_outs_valid : std_logic;
  signal extsi62_outs_ready : std_logic;
  signal source15_outs_valid : std_logic;
  signal source15_outs_ready : std_logic;
  signal constant54_outs : std_logic_vector(1 downto 0);
  signal constant54_outs_valid : std_logic;
  signal constant54_outs_ready : std_logic;
  signal extsi63_outs : std_logic_vector(5 downto 0);
  signal extsi63_outs_valid : std_logic;
  signal extsi63_outs_ready : std_logic;
  signal addi17_result : std_logic_vector(5 downto 0);
  signal addi17_result_valid : std_logic;
  signal addi17_result_ready : std_logic;
  signal buffer213_outs : std_logic_vector(5 downto 0);
  signal buffer213_outs_valid : std_logic;
  signal buffer213_outs_ready : std_logic;
  signal fork66_outs_0 : std_logic_vector(5 downto 0);
  signal fork66_outs_0_valid : std_logic;
  signal fork66_outs_0_ready : std_logic;
  signal fork66_outs_1 : std_logic_vector(5 downto 0);
  signal fork66_outs_1_valid : std_logic;
  signal fork66_outs_1_ready : std_logic;
  signal trunci21_outs : std_logic_vector(4 downto 0);
  signal trunci21_outs_valid : std_logic;
  signal trunci21_outs_ready : std_logic;
  signal cmpi4_result : std_logic_vector(0 downto 0);
  signal cmpi4_result_valid : std_logic;
  signal cmpi4_result_ready : std_logic;
  signal buffer214_outs : std_logic_vector(0 downto 0);
  signal buffer214_outs_valid : std_logic;
  signal buffer214_outs_ready : std_logic;
  signal fork67_outs_0 : std_logic_vector(0 downto 0);
  signal fork67_outs_0_valid : std_logic;
  signal fork67_outs_0_ready : std_logic;
  signal fork67_outs_1 : std_logic_vector(0 downto 0);
  signal fork67_outs_1_valid : std_logic;
  signal fork67_outs_1_ready : std_logic;
  signal fork67_outs_2 : std_logic_vector(0 downto 0);
  signal fork67_outs_2_valid : std_logic;
  signal fork67_outs_2_ready : std_logic;
  signal fork67_outs_3 : std_logic_vector(0 downto 0);
  signal fork67_outs_3_valid : std_logic;
  signal fork67_outs_3_ready : std_logic;
  signal fork67_outs_4 : std_logic_vector(0 downto 0);
  signal fork67_outs_4_valid : std_logic;
  signal fork67_outs_4_ready : std_logic;
  signal fork67_outs_5 : std_logic_vector(0 downto 0);
  signal fork67_outs_5_valid : std_logic;
  signal fork67_outs_5_ready : std_logic;
  signal fork67_outs_6 : std_logic_vector(0 downto 0);
  signal fork67_outs_6_valid : std_logic;
  signal fork67_outs_6_ready : std_logic;
  signal fork67_outs_7 : std_logic_vector(0 downto 0);
  signal fork67_outs_7_valid : std_logic;
  signal fork67_outs_7_ready : std_logic;
  signal cond_br27_trueOut : std_logic_vector(4 downto 0);
  signal cond_br27_trueOut_valid : std_logic;
  signal cond_br27_trueOut_ready : std_logic;
  signal cond_br27_falseOut : std_logic_vector(4 downto 0);
  signal cond_br27_falseOut_valid : std_logic;
  signal cond_br27_falseOut_ready : std_logic;
  signal buffer212_outs : std_logic_vector(31 downto 0);
  signal buffer212_outs_valid : std_logic;
  signal buffer212_outs_ready : std_logic;
  signal cond_br28_trueOut : std_logic_vector(31 downto 0);
  signal cond_br28_trueOut_valid : std_logic;
  signal cond_br28_trueOut_ready : std_logic;
  signal cond_br28_falseOut : std_logic_vector(31 downto 0);
  signal cond_br28_falseOut_valid : std_logic;
  signal cond_br28_falseOut_ready : std_logic;
  signal buffer174_outs : std_logic_vector(0 downto 0);
  signal buffer174_outs_valid : std_logic;
  signal buffer174_outs_ready : std_logic;
  signal cond_br29_trueOut : std_logic_vector(4 downto 0);
  signal cond_br29_trueOut_valid : std_logic;
  signal cond_br29_trueOut_ready : std_logic;
  signal cond_br29_falseOut : std_logic_vector(4 downto 0);
  signal cond_br29_falseOut_valid : std_logic;
  signal cond_br29_falseOut_ready : std_logic;
  signal cond_br30_trueOut_valid : std_logic;
  signal cond_br30_trueOut_ready : std_logic;
  signal cond_br30_falseOut_valid : std_logic;
  signal cond_br30_falseOut_ready : std_logic;
  signal buffer176_outs : std_logic_vector(0 downto 0);
  signal buffer176_outs_valid : std_logic;
  signal buffer176_outs_ready : std_logic;
  signal cond_br97_trueOut_valid : std_logic;
  signal cond_br97_trueOut_ready : std_logic;
  signal cond_br97_falseOut_valid : std_logic;
  signal cond_br97_falseOut_ready : std_logic;
  signal buffer177_outs : std_logic_vector(0 downto 0);
  signal buffer177_outs_valid : std_logic;
  signal buffer177_outs_ready : std_logic;
  signal cond_br98_trueOut_valid : std_logic;
  signal cond_br98_trueOut_ready : std_logic;
  signal cond_br98_falseOut_valid : std_logic;
  signal cond_br98_falseOut_ready : std_logic;
  signal cond_br99_trueOut_valid : std_logic;
  signal cond_br99_trueOut_ready : std_logic;
  signal cond_br99_falseOut_valid : std_logic;
  signal cond_br99_falseOut_ready : std_logic;
  signal extsi64_outs : std_logic_vector(5 downto 0);
  signal extsi64_outs_valid : std_logic;
  signal extsi64_outs_ready : std_logic;
  signal source16_outs_valid : std_logic;
  signal source16_outs_ready : std_logic;
  signal constant55_outs : std_logic_vector(4 downto 0);
  signal constant55_outs_valid : std_logic;
  signal constant55_outs_ready : std_logic;
  signal extsi65_outs : std_logic_vector(5 downto 0);
  signal extsi65_outs_valid : std_logic;
  signal extsi65_outs_ready : std_logic;
  signal source17_outs_valid : std_logic;
  signal source17_outs_ready : std_logic;
  signal constant56_outs : std_logic_vector(1 downto 0);
  signal constant56_outs_valid : std_logic;
  signal constant56_outs_ready : std_logic;
  signal extsi66_outs : std_logic_vector(5 downto 0);
  signal extsi66_outs_valid : std_logic;
  signal extsi66_outs_ready : std_logic;
  signal buffer216_outs : std_logic_vector(5 downto 0);
  signal buffer216_outs_valid : std_logic;
  signal buffer216_outs_ready : std_logic;
  signal addi18_result : std_logic_vector(5 downto 0);
  signal addi18_result_valid : std_logic;
  signal addi18_result_ready : std_logic;
  signal buffer217_outs : std_logic_vector(5 downto 0);
  signal buffer217_outs_valid : std_logic;
  signal buffer217_outs_ready : std_logic;
  signal fork68_outs_0 : std_logic_vector(5 downto 0);
  signal fork68_outs_0_valid : std_logic;
  signal fork68_outs_0_ready : std_logic;
  signal fork68_outs_1 : std_logic_vector(5 downto 0);
  signal fork68_outs_1_valid : std_logic;
  signal fork68_outs_1_ready : std_logic;
  signal trunci22_outs : std_logic_vector(4 downto 0);
  signal trunci22_outs_valid : std_logic;
  signal trunci22_outs_ready : std_logic;
  signal cmpi5_result : std_logic_vector(0 downto 0);
  signal cmpi5_result_valid : std_logic;
  signal cmpi5_result_ready : std_logic;
  signal buffer218_outs : std_logic_vector(0 downto 0);
  signal buffer218_outs_valid : std_logic;
  signal buffer218_outs_ready : std_logic;
  signal fork69_outs_0 : std_logic_vector(0 downto 0);
  signal fork69_outs_0_valid : std_logic;
  signal fork69_outs_0_ready : std_logic;
  signal fork69_outs_1 : std_logic_vector(0 downto 0);
  signal fork69_outs_1_valid : std_logic;
  signal fork69_outs_1_ready : std_logic;
  signal fork69_outs_2 : std_logic_vector(0 downto 0);
  signal fork69_outs_2_valid : std_logic;
  signal fork69_outs_2_ready : std_logic;
  signal fork69_outs_3 : std_logic_vector(0 downto 0);
  signal fork69_outs_3_valid : std_logic;
  signal fork69_outs_3_ready : std_logic;
  signal fork69_outs_4 : std_logic_vector(0 downto 0);
  signal fork69_outs_4_valid : std_logic;
  signal fork69_outs_4_ready : std_logic;
  signal fork69_outs_5 : std_logic_vector(0 downto 0);
  signal fork69_outs_5_valid : std_logic;
  signal fork69_outs_5_ready : std_logic;
  signal fork69_outs_6 : std_logic_vector(0 downto 0);
  signal fork69_outs_6_valid : std_logic;
  signal fork69_outs_6_ready : std_logic;
  signal cond_br31_trueOut : std_logic_vector(4 downto 0);
  signal cond_br31_trueOut_valid : std_logic;
  signal cond_br31_trueOut_ready : std_logic;
  signal cond_br31_falseOut : std_logic_vector(4 downto 0);
  signal cond_br31_falseOut_valid : std_logic;
  signal cond_br31_falseOut_ready : std_logic;
  signal cond_br32_trueOut : std_logic_vector(31 downto 0);
  signal cond_br32_trueOut_valid : std_logic;
  signal cond_br32_trueOut_ready : std_logic;
  signal cond_br32_falseOut : std_logic_vector(31 downto 0);
  signal cond_br32_falseOut_valid : std_logic;
  signal cond_br32_falseOut_ready : std_logic;
  signal cond_br33_trueOut_valid : std_logic;
  signal cond_br33_trueOut_ready : std_logic;
  signal cond_br33_falseOut_valid : std_logic;
  signal cond_br33_falseOut_ready : std_logic;
  signal buffer184_outs : std_logic_vector(0 downto 0);
  signal buffer184_outs_valid : std_logic;
  signal buffer184_outs_ready : std_logic;
  signal fork70_outs_0_valid : std_logic;
  signal fork70_outs_0_ready : std_logic;
  signal fork70_outs_1_valid : std_logic;
  signal fork70_outs_1_ready : std_logic;
  signal fork70_outs_2_valid : std_logic;
  signal fork70_outs_2_ready : std_logic;
  signal fork70_outs_3_valid : std_logic;
  signal fork70_outs_3_ready : std_logic;
  signal fork70_outs_4_valid : std_logic;
  signal fork70_outs_4_ready : std_logic;

begin

  tmp_end_valid <= mem_controller7_memEnd_valid;
  mem_controller7_memEnd_ready <= tmp_end_ready;
  A_end_valid <= mem_controller6_memEnd_valid;
  mem_controller6_memEnd_ready <= A_end_ready;
  B_end_valid <= mem_controller5_memEnd_valid;
  mem_controller5_memEnd_ready <= B_end_ready;
  C_end_valid <= mem_controller4_memEnd_valid;
  mem_controller4_memEnd_ready <= C_end_ready;
  D_end_valid <= mem_controller3_memEnd_valid;
  mem_controller3_memEnd_ready <= D_end_ready;
  end_valid <= fork0_outs_1_valid;
  fork0_outs_1_ready <= end_ready;
  tmp_loadEn <= mem_controller7_loadEn;
  tmp_loadAddr <= mem_controller7_loadAddr;
  tmp_storeEn <= mem_controller7_storeEn;
  tmp_storeAddr <= mem_controller7_storeAddr;
  tmp_storeData <= mem_controller7_storeData;
  A_loadEn <= mem_controller6_loadEn;
  A_loadAddr <= mem_controller6_loadAddr;
  A_storeEn <= mem_controller6_storeEn;
  A_storeAddr <= mem_controller6_storeAddr;
  A_storeData <= mem_controller6_storeData;
  B_loadEn <= mem_controller5_loadEn;
  B_loadAddr <= mem_controller5_loadAddr;
  B_storeEn <= mem_controller5_storeEn;
  B_storeAddr <= mem_controller5_storeAddr;
  B_storeData <= mem_controller5_storeData;
  C_loadEn <= mem_controller4_loadEn;
  C_loadAddr <= mem_controller4_loadAddr;
  C_storeEn <= mem_controller4_storeEn;
  C_storeAddr <= mem_controller4_storeAddr;
  C_storeData <= mem_controller4_storeData;
  D_loadEn <= mem_controller3_loadEn;
  D_loadAddr <= mem_controller3_loadAddr;
  D_storeEn <= mem_controller3_storeEn;
  D_storeAddr <= mem_controller3_storeAddr;
  D_storeData <= mem_controller3_storeData;

  fork0 : entity work.fork_dataless(arch) generic map(5)
    port map(
      ins_valid => start_valid,
      ins_ready => start_ready,
      clk => clk,
      rst => rst,
      outs_valid(0) => fork0_outs_0_valid,
      outs_valid(1) => fork0_outs_1_valid,
      outs_valid(2) => fork0_outs_2_valid,
      outs_valid(3) => fork0_outs_3_valid,
      outs_valid(4) => fork0_outs_4_valid,
      outs_ready(0) => fork0_outs_0_ready,
      outs_ready(1) => fork0_outs_1_ready,
      outs_ready(2) => fork0_outs_2_ready,
      outs_ready(3) => fork0_outs_3_ready,
      outs_ready(4) => fork0_outs_4_ready
    );

  mem_controller3 : entity work.mem_controller(arch) generic map(2, 2, 2, 32, 7)
    port map(
      loadData => D_loadData,
      memStart_valid => D_start_valid,
      memStart_ready => D_start_ready,
      ctrl(0) => extsi17_outs,
      ctrl(1) => extsi21_outs,
      ctrl_valid(0) => extsi17_outs_valid,
      ctrl_valid(1) => extsi21_outs_valid,
      ctrl_ready(0) => extsi17_outs_ready,
      ctrl_ready(1) => extsi21_outs_ready,
      ldAddr(0) => load3_addrOut,
      ldAddr(1) => load6_addrOut,
      ldAddr_valid(0) => load3_addrOut_valid,
      ldAddr_valid(1) => load6_addrOut_valid,
      ldAddr_ready(0) => load3_addrOut_ready,
      ldAddr_ready(1) => load6_addrOut_ready,
      stAddr(0) => store2_addrOut,
      stAddr(1) => store3_addrOut,
      stAddr_valid(0) => store2_addrOut_valid,
      stAddr_valid(1) => store3_addrOut_valid,
      stAddr_ready(0) => store2_addrOut_ready,
      stAddr_ready(1) => store3_addrOut_ready,
      stData(0) => store2_dataToMem,
      stData(1) => store3_dataToMem,
      stData_valid(0) => store2_dataToMem_valid,
      stData_valid(1) => store3_dataToMem_valid,
      stData_ready(0) => store2_dataToMem_ready,
      stData_ready(1) => store3_dataToMem_ready,
      ctrlEnd_valid => fork70_outs_4_valid,
      ctrlEnd_ready => fork70_outs_4_ready,
      clk => clk,
      rst => rst,
      ldData(0) => mem_controller3_ldData_0,
      ldData(1) => mem_controller3_ldData_1,
      ldData_valid(0) => mem_controller3_ldData_0_valid,
      ldData_valid(1) => mem_controller3_ldData_1_valid,
      ldData_ready(0) => mem_controller3_ldData_0_ready,
      ldData_ready(1) => mem_controller3_ldData_1_ready,
      stDone_valid(0) => mem_controller3_stDone_0_valid,
      stDone_valid(1) => mem_controller3_stDone_1_valid,
      stDone_ready(0) => mem_controller3_stDone_0_ready,
      stDone_ready(1) => mem_controller3_stDone_1_ready,
      memEnd_valid => mem_controller3_memEnd_valid,
      memEnd_ready => mem_controller3_memEnd_ready,
      loadEn => mem_controller3_loadEn,
      loadAddr => mem_controller3_loadAddr,
      storeEn => mem_controller3_storeEn,
      storeAddr => mem_controller3_storeAddr,
      storeData => mem_controller3_storeData
    );

  mem_controller4 : entity work.mem_controller_storeless(arch) generic map(1, 32, 7)
    port map(
      loadData => C_loadData,
      memStart_valid => C_start_valid,
      memStart_ready => C_start_ready,
      ldAddr(0) => load5_addrOut,
      ldAddr_valid(0) => load5_addrOut_valid,
      ldAddr_ready(0) => load5_addrOut_ready,
      ctrlEnd_valid => fork70_outs_3_valid,
      ctrlEnd_ready => fork70_outs_3_ready,
      clk => clk,
      rst => rst,
      ldData(0) => mem_controller4_ldData_0,
      ldData_valid(0) => mem_controller4_ldData_0_valid,
      ldData_ready(0) => mem_controller4_ldData_0_ready,
      memEnd_valid => mem_controller4_memEnd_valid,
      memEnd_ready => mem_controller4_memEnd_ready,
      loadEn => mem_controller4_loadEn,
      loadAddr => mem_controller4_loadAddr,
      storeEn => mem_controller4_storeEn,
      storeAddr => mem_controller4_storeAddr,
      storeData => mem_controller4_storeData
    );

  mem_controller5 : entity work.mem_controller_storeless(arch) generic map(1, 32, 7)
    port map(
      loadData => B_loadData,
      memStart_valid => B_start_valid,
      memStart_ready => B_start_ready,
      ldAddr(0) => load1_addrOut,
      ldAddr_valid(0) => load1_addrOut_valid,
      ldAddr_ready(0) => load1_addrOut_ready,
      ctrlEnd_valid => fork70_outs_2_valid,
      ctrlEnd_ready => fork70_outs_2_ready,
      clk => clk,
      rst => rst,
      ldData(0) => mem_controller5_ldData_0,
      ldData_valid(0) => mem_controller5_ldData_0_valid,
      ldData_ready(0) => mem_controller5_ldData_0_ready,
      memEnd_valid => mem_controller5_memEnd_valid,
      memEnd_ready => mem_controller5_memEnd_ready,
      loadEn => mem_controller5_loadEn,
      loadAddr => mem_controller5_loadAddr,
      storeEn => mem_controller5_storeEn,
      storeAddr => mem_controller5_storeAddr,
      storeData => mem_controller5_storeData
    );

  mem_controller6 : entity work.mem_controller_storeless(arch) generic map(1, 32, 7)
    port map(
      loadData => A_loadData,
      memStart_valid => A_start_valid,
      memStart_ready => A_start_ready,
      ldAddr(0) => load0_addrOut,
      ldAddr_valid(0) => load0_addrOut_valid,
      ldAddr_ready(0) => load0_addrOut_ready,
      ctrlEnd_valid => fork70_outs_1_valid,
      ctrlEnd_ready => fork70_outs_1_ready,
      clk => clk,
      rst => rst,
      ldData(0) => mem_controller6_ldData_0,
      ldData_valid(0) => mem_controller6_ldData_0_valid,
      ldData_ready(0) => mem_controller6_ldData_0_ready,
      memEnd_valid => mem_controller6_memEnd_valid,
      memEnd_ready => mem_controller6_memEnd_ready,
      loadEn => mem_controller6_loadEn,
      loadAddr => mem_controller6_loadAddr,
      storeEn => mem_controller6_storeEn,
      storeAddr => mem_controller6_storeAddr,
      storeData => mem_controller6_storeData
    );

  mem_controller7 : entity work.mem_controller(arch) generic map(2, 2, 2, 32, 7)
    port map(
      loadData => tmp_loadData,
      memStart_valid => tmp_start_valid,
      memStart_ready => tmp_start_ready,
      ctrl(0) => extsi2_outs,
      ctrl(1) => extsi7_outs,
      ctrl_valid(0) => extsi2_outs_valid,
      ctrl_valid(1) => extsi7_outs_valid,
      ctrl_ready(0) => extsi2_outs_ready,
      ctrl_ready(1) => extsi7_outs_ready,
      stAddr(0) => store0_addrOut,
      stAddr(1) => store1_addrOut,
      stAddr_valid(0) => store0_addrOut_valid,
      stAddr_valid(1) => store1_addrOut_valid,
      stAddr_ready(0) => store0_addrOut_ready,
      stAddr_ready(1) => store1_addrOut_ready,
      stData(0) => store0_dataToMem,
      stData(1) => store1_dataToMem,
      stData_valid(0) => store0_dataToMem_valid,
      stData_valid(1) => store1_dataToMem_valid,
      stData_ready(0) => store0_dataToMem_ready,
      stData_ready(1) => store1_dataToMem_ready,
      ldAddr(0) => load2_addrOut,
      ldAddr(1) => load4_addrOut,
      ldAddr_valid(0) => load2_addrOut_valid,
      ldAddr_valid(1) => load4_addrOut_valid,
      ldAddr_ready(0) => load2_addrOut_ready,
      ldAddr_ready(1) => load4_addrOut_ready,
      ctrlEnd_valid => fork70_outs_0_valid,
      ctrlEnd_ready => fork70_outs_0_ready,
      clk => clk,
      rst => rst,
      stDone_valid(0) => mem_controller7_stDone_0_valid,
      stDone_valid(1) => mem_controller7_stDone_1_valid,
      stDone_ready(0) => mem_controller7_stDone_0_ready,
      stDone_ready(1) => mem_controller7_stDone_1_ready,
      ldData(0) => mem_controller7_ldData_0,
      ldData(1) => mem_controller7_ldData_1,
      ldData_valid(0) => mem_controller7_ldData_0_valid,
      ldData_valid(1) => mem_controller7_ldData_1_valid,
      ldData_ready(0) => mem_controller7_ldData_0_ready,
      ldData_ready(1) => mem_controller7_ldData_1_ready,
      memEnd_valid => mem_controller7_memEnd_valid,
      memEnd_ready => mem_controller7_memEnd_ready,
      loadEn => mem_controller7_loadEn,
      loadAddr => mem_controller7_loadAddr,
      storeEn => mem_controller7_storeEn,
      storeAddr => mem_controller7_storeAddr,
      storeData => mem_controller7_storeData
    );

  constant29 : entity work.handshake_constant_0(arch) generic map(1)
    port map(
      ctrl_valid => fork0_outs_0_valid,
      ctrl_ready => fork0_outs_0_ready,
      clk => clk,
      rst => rst,
      outs => constant29_outs,
      outs_valid => constant29_outs_valid,
      outs_ready => constant29_outs_ready
    );

  extsi34 : entity work.extsi(arch) generic map(1, 5)
    port map(
      ins => constant29_outs,
      ins_valid => constant29_outs_valid,
      ins_ready => constant29_outs_ready,
      clk => clk,
      rst => rst,
      outs => extsi34_outs,
      outs_valid => extsi34_outs_valid,
      outs_ready => extsi34_outs_ready
    );

  mux25 : entity work.mux_dataless(arch) generic map(2, 1)
    port map(
      index => init0_outs,
      index_valid => init0_outs_valid,
      index_ready => init0_outs_ready,
      ins_valid(0) => fork0_outs_3_valid,
      ins_valid(1) => cond_br88_trueOut_valid,
      ins_ready(0) => fork0_outs_3_ready,
      ins_ready(1) => cond_br88_trueOut_ready,
      clk => clk,
      rst => rst,
      outs_valid => mux25_outs_valid,
      outs_ready => mux25_outs_ready
    );

  init0 : entity work.tehb_init(arch) generic map(1, 0)
    port map(
      ins => fork30_outs_3,
      ins_valid => fork30_outs_3_valid,
      ins_ready => fork30_outs_3_ready,
      clk => clk,
      rst => rst,
      outs => init0_outs,
      outs_valid => init0_outs_valid,
      outs_ready => init0_outs_ready
    );

  mux0 : entity work.mux(arch) generic map(2, 5, 1)
    port map(
      index => fork1_outs_0,
      index_valid => fork1_outs_0_valid,
      index_ready => fork1_outs_0_ready,
      ins(0) => extsi34_outs,
      ins(1) => cond_br17_trueOut,
      ins_valid(0) => extsi34_outs_valid,
      ins_valid(1) => cond_br17_trueOut_valid,
      ins_ready(0) => extsi34_outs_ready,
      ins_ready(1) => cond_br17_trueOut_ready,
      clk => clk,
      rst => rst,
      outs => mux0_outs,
      outs_valid => mux0_outs_valid,
      outs_ready => mux0_outs_ready
    );

  mux1 : entity work.mux(arch) generic map(2, 32, 1)
    port map(
      index => buffer7_outs,
      index_valid => buffer7_outs_valid,
      index_ready => buffer7_outs_ready,
      ins(0) => alpha,
      ins(1) => cond_br18_trueOut,
      ins_valid(0) => alpha_valid,
      ins_valid(1) => cond_br18_trueOut_valid,
      ins_ready(0) => alpha_ready,
      ins_ready(1) => cond_br18_trueOut_ready,
      clk => clk,
      rst => rst,
      outs => mux1_outs,
      outs_valid => mux1_outs_valid,
      outs_ready => mux1_outs_ready
    );

  buffer7 : entity work.tfifo(arch) generic map(1, 1)
    port map(
      ins => fork1_outs_1,
      ins_valid => fork1_outs_1_valid,
      ins_ready => fork1_outs_1_ready,
      clk => clk,
      rst => rst,
      outs => buffer7_outs,
      outs_valid => buffer7_outs_valid,
      outs_ready => buffer7_outs_ready
    );

  mux2 : entity work.mux(arch) generic map(2, 32, 1)
    port map(
      index => buffer8_outs,
      index_valid => buffer8_outs_valid,
      index_ready => buffer8_outs_ready,
      ins(0) => beta,
      ins(1) => cond_br19_trueOut,
      ins_valid(0) => beta_valid,
      ins_valid(1) => cond_br19_trueOut_valid,
      ins_ready(0) => beta_ready,
      ins_ready(1) => cond_br19_trueOut_ready,
      clk => clk,
      rst => rst,
      outs => mux2_outs,
      outs_valid => mux2_outs_valid,
      outs_ready => mux2_outs_ready
    );

  buffer8 : entity work.tfifo(arch) generic map(1, 1)
    port map(
      ins => fork1_outs_2,
      ins_valid => fork1_outs_2_valid,
      ins_ready => fork1_outs_2_ready,
      clk => clk,
      rst => rst,
      outs => buffer8_outs,
      outs_valid => buffer8_outs_valid,
      outs_ready => buffer8_outs_ready
    );

  control_merge0 : entity work.control_merge_dataless(arch) generic map(2, 1)
    port map(
      ins_valid(0) => fork0_outs_4_valid,
      ins_valid(1) => cond_br20_trueOut_valid,
      ins_ready(0) => fork0_outs_4_ready,
      ins_ready(1) => cond_br20_trueOut_ready,
      clk => clk,
      rst => rst,
      outs_valid => control_merge0_outs_valid,
      outs_ready => control_merge0_outs_ready,
      index => control_merge0_index,
      index_valid => control_merge0_index_valid,
      index_ready => control_merge0_index_ready
    );

  fork1 : entity work.handshake_fork(arch) generic map(3, 1)
    port map(
      ins => control_merge0_index,
      ins_valid => control_merge0_index_valid,
      ins_ready => control_merge0_index_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork1_outs_0,
      outs(1) => fork1_outs_1,
      outs(2) => fork1_outs_2,
      outs_valid(0) => fork1_outs_0_valid,
      outs_valid(1) => fork1_outs_1_valid,
      outs_valid(2) => fork1_outs_2_valid,
      outs_ready(0) => fork1_outs_0_ready,
      outs_ready(1) => fork1_outs_1_ready,
      outs_ready(2) => fork1_outs_2_ready
    );

  fork2 : entity work.fork_dataless(arch) generic map(2)
    port map(
      ins_valid => control_merge0_outs_valid,
      ins_ready => control_merge0_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid(0) => fork2_outs_0_valid,
      outs_valid(1) => fork2_outs_1_valid,
      outs_ready(0) => fork2_outs_0_ready,
      outs_ready(1) => fork2_outs_1_ready
    );

  constant30 : entity work.handshake_constant_0(arch) generic map(1)
    port map(
      ctrl_valid => fork2_outs_0_valid,
      ctrl_ready => fork2_outs_0_ready,
      clk => clk,
      rst => rst,
      outs => constant30_outs,
      outs_valid => constant30_outs_valid,
      outs_ready => constant30_outs_ready
    );

  extsi33 : entity work.extsi(arch) generic map(1, 5)
    port map(
      ins => constant30_outs,
      ins_valid => constant30_outs_valid,
      ins_ready => constant30_outs_ready,
      clk => clk,
      rst => rst,
      outs => extsi33_outs,
      outs_valid => extsi33_outs_valid,
      outs_ready => extsi33_outs_ready
    );

  buffer10 : entity work.tehb(arch) generic map(32)
    port map(
      ins => mux1_outs,
      ins_valid => mux1_outs_valid,
      ins_ready => mux1_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer10_outs,
      outs_valid => buffer10_outs_valid,
      outs_ready => buffer10_outs_ready
    );

  buffer11 : entity work.oehb(arch) generic map(32)
    port map(
      ins => mux2_outs,
      ins_valid => mux2_outs_valid,
      ins_ready => mux2_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer11_outs,
      outs_valid => buffer11_outs_valid,
      outs_ready => buffer11_outs_ready
    );

  buffer14 : entity work.tehb(arch) generic map(32)
    port map(
      ins => buffer11_outs,
      ins_valid => buffer11_outs_valid,
      ins_ready => buffer11_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer14_outs,
      outs_valid => buffer14_outs_valid,
      outs_ready => buffer14_outs_ready
    );

  buffer6 : entity work.tehb(arch) generic map(5)
    port map(
      ins => mux0_outs,
      ins_valid => mux0_outs_valid,
      ins_ready => mux0_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer6_outs,
      outs_valid => buffer6_outs_valid,
      outs_ready => buffer6_outs_ready
    );

  buffer5 : entity work.tehb_dataless(arch)
    port map(
      ins_valid => mux25_outs_valid,
      ins_ready => mux25_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer5_outs_valid,
      outs_ready => buffer5_outs_ready
    );

  mux30 : entity work.mux_dataless(arch) generic map(2, 1)
    port map(
      index => init5_outs,
      index_valid => init5_outs_valid,
      index_ready => init5_outs_ready,
      ins_valid(0) => buffer5_outs_valid,
      ins_valid(1) => cond_br85_trueOut_valid,
      ins_ready(0) => buffer5_outs_ready,
      ins_ready(1) => cond_br85_trueOut_ready,
      clk => clk,
      rst => rst,
      outs_valid => mux30_outs_valid,
      outs_ready => mux30_outs_ready
    );

  init5 : entity work.tehb_init(arch) generic map(1, 0)
    port map(
      ins => buffer9_outs,
      ins_valid => buffer9_outs_valid,
      ins_ready => buffer9_outs_ready,
      clk => clk,
      rst => rst,
      outs => init5_outs,
      outs_valid => init5_outs_valid,
      outs_ready => init5_outs_ready
    );

  buffer9 : entity work.tfifo(arch) generic map(1, 1)
    port map(
      ins => fork27_outs_4,
      ins_valid => fork27_outs_4_valid,
      ins_ready => fork27_outs_4_ready,
      clk => clk,
      rst => rst,
      outs => buffer9_outs,
      outs_valid => buffer9_outs_valid,
      outs_ready => buffer9_outs_ready
    );

  mux3 : entity work.mux(arch) generic map(2, 5, 1)
    port map(
      index => fork6_outs_1,
      index_valid => fork6_outs_1_valid,
      index_ready => fork6_outs_1_ready,
      ins(0) => extsi33_outs,
      ins(1) => cond_br12_trueOut,
      ins_valid(0) => extsi33_outs_valid,
      ins_valid(1) => cond_br12_trueOut_valid,
      ins_ready(0) => extsi33_outs_ready,
      ins_ready(1) => cond_br12_trueOut_ready,
      clk => clk,
      rst => rst,
      outs => mux3_outs,
      outs_valid => mux3_outs_valid,
      outs_ready => mux3_outs_ready
    );

  buffer18 : entity work.tehb(arch) generic map(5)
    port map(
      ins => mux3_outs,
      ins_valid => mux3_outs_valid,
      ins_ready => mux3_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer18_outs,
      outs_valid => buffer18_outs_valid,
      outs_ready => buffer18_outs_ready
    );

  fork3 : entity work.handshake_fork(arch) generic map(2, 5)
    port map(
      ins => buffer18_outs,
      ins_valid => buffer18_outs_valid,
      ins_ready => buffer18_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork3_outs_0,
      outs(1) => fork3_outs_1,
      outs_valid(0) => fork3_outs_0_valid,
      outs_valid(1) => fork3_outs_1_valid,
      outs_ready(0) => fork3_outs_0_ready,
      outs_ready(1) => fork3_outs_1_ready
    );

  extsi35 : entity work.extsi(arch) generic map(5, 7)
    port map(
      ins => fork3_outs_0,
      ins_valid => fork3_outs_0_valid,
      ins_ready => fork3_outs_0_ready,
      clk => clk,
      rst => rst,
      outs => extsi35_outs,
      outs_valid => extsi35_outs_valid,
      outs_ready => extsi35_outs_ready
    );

  buffer15 : entity work.oehb(arch) generic map(32)
    port map(
      ins => buffer10_outs,
      ins_valid => buffer10_outs_valid,
      ins_ready => buffer10_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer15_outs,
      outs_valid => buffer15_outs_valid,
      outs_ready => buffer15_outs_ready
    );

  mux4 : entity work.mux(arch) generic map(2, 32, 1)
    port map(
      index => buffer12_outs,
      index_valid => buffer12_outs_valid,
      index_ready => buffer12_outs_ready,
      ins(0) => buffer15_outs,
      ins(1) => cond_br13_trueOut,
      ins_valid(0) => buffer15_outs_valid,
      ins_valid(1) => cond_br13_trueOut_valid,
      ins_ready(0) => buffer15_outs_ready,
      ins_ready(1) => cond_br13_trueOut_ready,
      clk => clk,
      rst => rst,
      outs => mux4_outs,
      outs_valid => mux4_outs_valid,
      outs_ready => mux4_outs_ready
    );

  buffer12 : entity work.tfifo(arch) generic map(1, 1)
    port map(
      ins => fork6_outs_2,
      ins_valid => fork6_outs_2_valid,
      ins_ready => fork6_outs_2_ready,
      clk => clk,
      rst => rst,
      outs => buffer12_outs,
      outs_valid => buffer12_outs_valid,
      outs_ready => buffer12_outs_ready
    );

  mux5 : entity work.mux(arch) generic map(2, 32, 1)
    port map(
      index => buffer13_outs,
      index_valid => buffer13_outs_valid,
      index_ready => buffer13_outs_ready,
      ins(0) => buffer14_outs,
      ins(1) => cond_br14_trueOut,
      ins_valid(0) => buffer14_outs_valid,
      ins_valid(1) => cond_br14_trueOut_valid,
      ins_ready(0) => buffer14_outs_ready,
      ins_ready(1) => cond_br14_trueOut_ready,
      clk => clk,
      rst => rst,
      outs => mux5_outs,
      outs_valid => mux5_outs_valid,
      outs_ready => mux5_outs_ready
    );

  buffer13 : entity work.tfifo(arch) generic map(1, 1)
    port map(
      ins => fork6_outs_3,
      ins_valid => fork6_outs_3_valid,
      ins_ready => fork6_outs_3_ready,
      clk => clk,
      rst => rst,
      outs => buffer13_outs,
      outs_valid => buffer13_outs_valid,
      outs_ready => buffer13_outs_ready
    );

  mux6 : entity work.mux(arch) generic map(2, 5, 1)
    port map(
      index => fork6_outs_0,
      index_valid => fork6_outs_0_valid,
      index_ready => fork6_outs_0_ready,
      ins(0) => buffer6_outs,
      ins(1) => cond_br15_trueOut,
      ins_valid(0) => buffer6_outs_valid,
      ins_valid(1) => cond_br15_trueOut_valid,
      ins_ready(0) => buffer6_outs_ready,
      ins_ready(1) => cond_br15_trueOut_ready,
      clk => clk,
      rst => rst,
      outs => mux6_outs,
      outs_valid => mux6_outs_valid,
      outs_ready => mux6_outs_ready
    );

  buffer21 : entity work.oehb(arch) generic map(5)
    port map(
      ins => mux6_outs,
      ins_valid => mux6_outs_valid,
      ins_ready => mux6_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer21_outs,
      outs_valid => buffer21_outs_valid,
      outs_ready => buffer21_outs_ready
    );

  buffer24 : entity work.tehb(arch) generic map(5)
    port map(
      ins => buffer21_outs,
      ins_valid => buffer21_outs_valid,
      ins_ready => buffer21_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer24_outs,
      outs_valid => buffer24_outs_valid,
      outs_ready => buffer24_outs_ready
    );

  fork4 : entity work.handshake_fork(arch) generic map(2, 5)
    port map(
      ins => buffer24_outs,
      ins_valid => buffer24_outs_valid,
      ins_ready => buffer24_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork4_outs_0,
      outs(1) => fork4_outs_1,
      outs_valid(0) => fork4_outs_0_valid,
      outs_valid(1) => fork4_outs_1_valid,
      outs_ready(0) => fork4_outs_0_ready,
      outs_ready(1) => fork4_outs_1_ready
    );

  extsi36 : entity work.extsi(arch) generic map(5, 32)
    port map(
      ins => fork4_outs_1,
      ins_valid => fork4_outs_1_valid,
      ins_ready => fork4_outs_1_ready,
      clk => clk,
      rst => rst,
      outs => extsi36_outs,
      outs_valid => extsi36_outs_valid,
      outs_ready => extsi36_outs_ready
    );

  fork5 : entity work.handshake_fork(arch) generic map(2, 32)
    port map(
      ins => extsi36_outs,
      ins_valid => extsi36_outs_valid,
      ins_ready => extsi36_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork5_outs_0,
      outs(1) => fork5_outs_1,
      outs_valid(0) => fork5_outs_0_valid,
      outs_valid(1) => fork5_outs_1_valid,
      outs_ready(0) => fork5_outs_0_ready,
      outs_ready(1) => fork5_outs_1_ready
    );

  control_merge1 : entity work.control_merge_dataless(arch) generic map(2, 1)
    port map(
      ins_valid(0) => fork2_outs_1_valid,
      ins_valid(1) => cond_br16_trueOut_valid,
      ins_ready(0) => fork2_outs_1_ready,
      ins_ready(1) => cond_br16_trueOut_ready,
      clk => clk,
      rst => rst,
      outs_valid => control_merge1_outs_valid,
      outs_ready => control_merge1_outs_ready,
      index => control_merge1_index,
      index_valid => control_merge1_index_valid,
      index_ready => control_merge1_index_ready
    );

  fork6 : entity work.handshake_fork(arch) generic map(4, 1)
    port map(
      ins => control_merge1_index,
      ins_valid => control_merge1_index_valid,
      ins_ready => control_merge1_index_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork6_outs_0,
      outs(1) => fork6_outs_1,
      outs(2) => fork6_outs_2,
      outs(3) => fork6_outs_3,
      outs_valid(0) => fork6_outs_0_valid,
      outs_valid(1) => fork6_outs_1_valid,
      outs_valid(2) => fork6_outs_2_valid,
      outs_valid(3) => fork6_outs_3_valid,
      outs_ready(0) => fork6_outs_0_ready,
      outs_ready(1) => fork6_outs_1_ready,
      outs_ready(2) => fork6_outs_2_ready,
      outs_ready(3) => fork6_outs_3_ready
    );

  fork7 : entity work.fork_dataless(arch) generic map(3)
    port map(
      ins_valid => control_merge1_outs_valid,
      ins_ready => control_merge1_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid(0) => fork7_outs_0_valid,
      outs_valid(1) => fork7_outs_1_valid,
      outs_valid(2) => fork7_outs_2_valid,
      outs_ready(0) => fork7_outs_0_ready,
      outs_ready(1) => fork7_outs_1_ready,
      outs_ready(2) => fork7_outs_2_ready
    );

  constant31 : entity work.handshake_constant_1(arch) generic map(2)
    port map(
      ctrl_valid => fork7_outs_1_valid,
      ctrl_ready => fork7_outs_1_ready,
      clk => clk,
      rst => rst,
      outs => constant31_outs,
      outs_valid => constant31_outs_valid,
      outs_ready => constant31_outs_ready
    );

  extsi2 : entity work.extsi(arch) generic map(2, 32)
    port map(
      ins => constant31_outs,
      ins_valid => constant31_outs_valid,
      ins_ready => constant31_outs_ready,
      clk => clk,
      rst => rst,
      outs => extsi2_outs,
      outs_valid => extsi2_outs_valid,
      outs_ready => extsi2_outs_ready
    );

  constant32 : entity work.handshake_constant_0(arch) generic map(1)
    port map(
      ctrl_valid => fork7_outs_0_valid,
      ctrl_ready => fork7_outs_0_ready,
      clk => clk,
      rst => rst,
      outs => constant32_outs,
      outs_valid => constant32_outs_valid,
      outs_ready => constant32_outs_ready
    );

  fork8 : entity work.handshake_fork(arch) generic map(2, 1)
    port map(
      ins => constant32_outs,
      ins_valid => constant32_outs_valid,
      ins_ready => constant32_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork8_outs_0,
      outs(1) => fork8_outs_1,
      outs_valid(0) => fork8_outs_0_valid,
      outs_valid(1) => fork8_outs_1_valid,
      outs_ready(0) => fork8_outs_0_ready,
      outs_ready(1) => fork8_outs_1_ready
    );

  extsi4 : entity work.extsi(arch) generic map(1, 32)
    port map(
      ins => fork8_outs_1,
      ins_valid => fork8_outs_1_valid,
      ins_ready => fork8_outs_1_ready,
      clk => clk,
      rst => rst,
      outs => extsi4_outs,
      outs_valid => extsi4_outs_valid,
      outs_ready => extsi4_outs_ready
    );

  source0 : entity work.source(arch)
    port map(
      clk => clk,
      rst => rst,
      outs_valid => source0_outs_valid,
      outs_ready => source0_outs_ready
    );

  constant33 : entity work.handshake_constant_1(arch) generic map(2)
    port map(
      ctrl_valid => source0_outs_valid,
      ctrl_ready => source0_outs_ready,
      clk => clk,
      rst => rst,
      outs => constant33_outs,
      outs_valid => constant33_outs_valid,
      outs_ready => constant33_outs_ready
    );

  extsi5 : entity work.extsi(arch) generic map(2, 32)
    port map(
      ins => constant33_outs,
      ins_valid => constant33_outs_valid,
      ins_ready => constant33_outs_ready,
      clk => clk,
      rst => rst,
      outs => extsi5_outs,
      outs_valid => extsi5_outs_valid,
      outs_ready => extsi5_outs_ready
    );

  source1 : entity work.source(arch)
    port map(
      clk => clk,
      rst => rst,
      outs_valid => source1_outs_valid,
      outs_ready => source1_outs_ready
    );

  constant34 : entity work.handshake_constant_2(arch) generic map(3)
    port map(
      ctrl_valid => source1_outs_valid,
      ctrl_ready => source1_outs_ready,
      clk => clk,
      rst => rst,
      outs => constant34_outs,
      outs_valid => constant34_outs_valid,
      outs_ready => constant34_outs_ready
    );

  extsi6 : entity work.extsi(arch) generic map(3, 32)
    port map(
      ins => constant34_outs,
      ins_valid => constant34_outs_valid,
      ins_ready => constant34_outs_ready,
      clk => clk,
      rst => rst,
      outs => extsi6_outs,
      outs_valid => extsi6_outs_valid,
      outs_ready => extsi6_outs_ready
    );

  shli0 : entity work.shli(arch) generic map(32)
    port map(
      lhs => fork5_outs_0,
      lhs_valid => fork5_outs_0_valid,
      lhs_ready => fork5_outs_0_ready,
      rhs => extsi5_outs,
      rhs_valid => extsi5_outs_valid,
      rhs_ready => extsi5_outs_ready,
      clk => clk,
      rst => rst,
      result => shli0_result,
      result_valid => shli0_result_valid,
      result_ready => shli0_result_ready
    );

  buffer27 : entity work.oehb(arch) generic map(32)
    port map(
      ins => shli0_result,
      ins_valid => shli0_result_valid,
      ins_ready => shli0_result_ready,
      clk => clk,
      rst => rst,
      outs => buffer27_outs,
      outs_valid => buffer27_outs_valid,
      outs_ready => buffer27_outs_ready
    );

  trunci0 : entity work.trunci(arch) generic map(32, 7)
    port map(
      ins => buffer27_outs,
      ins_valid => buffer27_outs_valid,
      ins_ready => buffer27_outs_ready,
      clk => clk,
      rst => rst,
      outs => trunci0_outs,
      outs_valid => trunci0_outs_valid,
      outs_ready => trunci0_outs_ready
    );

  shli1 : entity work.shli(arch) generic map(32)
    port map(
      lhs => fork5_outs_1,
      lhs_valid => fork5_outs_1_valid,
      lhs_ready => fork5_outs_1_ready,
      rhs => extsi6_outs,
      rhs_valid => extsi6_outs_valid,
      rhs_ready => extsi6_outs_ready,
      clk => clk,
      rst => rst,
      result => shli1_result,
      result_valid => shli1_result_valid,
      result_ready => shli1_result_ready
    );

  buffer29 : entity work.oehb(arch) generic map(32)
    port map(
      ins => shli1_result,
      ins_valid => shli1_result_valid,
      ins_ready => shli1_result_ready,
      clk => clk,
      rst => rst,
      outs => buffer29_outs,
      outs_valid => buffer29_outs_valid,
      outs_ready => buffer29_outs_ready
    );

  trunci1 : entity work.trunci(arch) generic map(32, 7)
    port map(
      ins => buffer29_outs,
      ins_valid => buffer29_outs_valid,
      ins_ready => buffer29_outs_ready,
      clk => clk,
      rst => rst,
      outs => trunci1_outs,
      outs_valid => trunci1_outs_valid,
      outs_ready => trunci1_outs_ready
    );

  addi19 : entity work.addi(arch) generic map(7)
    port map(
      lhs => trunci0_outs,
      lhs_valid => trunci0_outs_valid,
      lhs_ready => trunci0_outs_ready,
      rhs => trunci1_outs,
      rhs_valid => trunci1_outs_valid,
      rhs_ready => trunci1_outs_ready,
      clk => clk,
      rst => rst,
      result => addi19_result,
      result_valid => addi19_result_valid,
      result_ready => addi19_result_ready
    );

  buffer30 : entity work.oehb(arch) generic map(7)
    port map(
      ins => addi19_result,
      ins_valid => addi19_result_valid,
      ins_ready => addi19_result_ready,
      clk => clk,
      rst => rst,
      outs => buffer30_outs,
      outs_valid => buffer30_outs_valid,
      outs_ready => buffer30_outs_ready
    );

  addi2 : entity work.addi(arch) generic map(7)
    port map(
      lhs => extsi35_outs,
      lhs_valid => extsi35_outs_valid,
      lhs_ready => extsi35_outs_ready,
      rhs => buffer30_outs,
      rhs_valid => buffer30_outs_valid,
      rhs_ready => buffer30_outs_ready,
      clk => clk,
      rst => rst,
      result => addi2_result,
      result_valid => addi2_result_valid,
      result_ready => addi2_result_ready
    );

  buffer0 : entity work.tfifo_dataless(arch) generic map(1)
    port map(
      ins_valid => store0_doneOut_valid,
      ins_ready => store0_doneOut_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer0_outs_valid,
      outs_ready => buffer0_outs_ready
    );

  fork9 : entity work.fork_dataless(arch) generic map(2)
    port map(
      ins_valid => buffer0_outs_valid,
      ins_ready => buffer0_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid(0) => fork9_outs_0_valid,
      outs_valid(1) => fork9_outs_1_valid,
      outs_ready(0) => fork9_outs_0_ready,
      outs_ready(1) => fork9_outs_1_ready
    );

  buffer31 : entity work.oehb(arch) generic map(7)
    port map(
      ins => addi2_result,
      ins_valid => addi2_result_valid,
      ins_ready => addi2_result_ready,
      clk => clk,
      rst => rst,
      outs => buffer31_outs,
      outs_valid => buffer31_outs_valid,
      outs_ready => buffer31_outs_ready
    );

  store0 : entity work.store(arch) generic map(32, 7)
    port map(
      addrIn => buffer31_outs,
      addrIn_valid => buffer31_outs_valid,
      addrIn_ready => buffer31_outs_ready,
      dataIn => extsi4_outs,
      dataIn_valid => extsi4_outs_valid,
      dataIn_ready => extsi4_outs_ready,
      doneFromMem_valid => mem_controller7_stDone_0_valid,
      doneFromMem_ready => mem_controller7_stDone_0_ready,
      clk => clk,
      rst => rst,
      addrOut => store0_addrOut,
      addrOut_valid => store0_addrOut_valid,
      addrOut_ready => store0_addrOut_ready,
      dataToMem => store0_dataToMem,
      dataToMem_valid => store0_dataToMem_valid,
      dataToMem_ready => store0_dataToMem_ready,
      doneOut_valid => store0_doneOut_valid,
      doneOut_ready => store0_doneOut_ready
    );

  extsi32 : entity work.extsi(arch) generic map(1, 5)
    port map(
      ins => fork8_outs_0,
      ins_valid => fork8_outs_0_valid,
      ins_ready => fork8_outs_0_ready,
      clk => clk,
      rst => rst,
      outs => extsi32_outs,
      outs_valid => extsi32_outs_valid,
      outs_ready => extsi32_outs_ready
    );

  buffer19 : entity work.tehb(arch) generic map(32)
    port map(
      ins => mux4_outs,
      ins_valid => mux4_outs_valid,
      ins_ready => mux4_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer19_outs,
      outs_valid => buffer19_outs_valid,
      outs_ready => buffer19_outs_ready
    );

  buffer20 : entity work.tehb(arch) generic map(32)
    port map(
      ins => mux5_outs,
      ins_valid => mux5_outs_valid,
      ins_ready => mux5_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer20_outs,
      outs_valid => buffer20_outs_valid,
      outs_ready => buffer20_outs_ready
    );

  cond_br83 : entity work.cond_br_dataless(arch)
    port map(
      condition => buffer22_outs,
      condition_valid => buffer22_outs_valid,
      condition_ready => buffer22_outs_ready,
      data_valid => fork11_outs_2_valid,
      data_ready => fork11_outs_2_ready,
      clk => clk,
      rst => rst,
      trueOut_valid => cond_br83_trueOut_valid,
      trueOut_ready => cond_br83_trueOut_ready,
      falseOut_valid => cond_br83_falseOut_valid,
      falseOut_ready => cond_br83_falseOut_ready
    );

  buffer22 : entity work.tfifo(arch) generic map(5, 1)
    port map(
      ins => fork25_outs_5,
      ins_valid => fork25_outs_5_valid,
      ins_ready => fork25_outs_5_ready,
      clk => clk,
      rst => rst,
      outs => buffer22_outs,
      outs_valid => buffer22_outs_valid,
      outs_ready => buffer22_outs_ready
    );

  sink0 : entity work.sink_dataless(arch)
    port map(
      ins_valid => cond_br83_falseOut_valid,
      ins_ready => cond_br83_falseOut_ready,
      clk => clk,
      rst => rst
    );

  buffer100 : entity work.oehb_dataless(arch)
    port map(
      ins_valid => buffer1_outs_valid,
      ins_ready => buffer1_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer100_outs_valid,
      outs_ready => buffer100_outs_ready
    );

  cond_br84 : entity work.cond_br_dataless(arch)
    port map(
      condition => buffer23_outs,
      condition_valid => buffer23_outs_valid,
      condition_ready => buffer23_outs_ready,
      data_valid => buffer100_outs_valid,
      data_ready => buffer100_outs_ready,
      clk => clk,
      rst => rst,
      trueOut_valid => cond_br84_trueOut_valid,
      trueOut_ready => cond_br84_trueOut_ready,
      falseOut_valid => cond_br84_falseOut_valid,
      falseOut_ready => cond_br84_falseOut_ready
    );

  buffer23 : entity work.tfifo(arch) generic map(5, 1)
    port map(
      ins => fork25_outs_4,
      ins_valid => fork25_outs_4_valid,
      ins_ready => fork25_outs_4_ready,
      clk => clk,
      rst => rst,
      outs => buffer23_outs,
      outs_valid => buffer23_outs_valid,
      outs_ready => buffer23_outs_ready
    );

  init10 : entity work.tehb_init(arch) generic map(1, 0)
    port map(
      ins => fork25_outs_3,
      ins_valid => fork25_outs_3_valid,
      ins_ready => fork25_outs_3_ready,
      clk => clk,
      rst => rst,
      outs => init10_outs,
      outs_valid => init10_outs_valid,
      outs_ready => init10_outs_ready
    );

  fork10 : entity work.handshake_fork(arch) generic map(2, 1)
    port map(
      ins => init10_outs,
      ins_valid => init10_outs_valid,
      ins_ready => init10_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork10_outs_0,
      outs(1) => fork10_outs_1,
      outs_valid(0) => fork10_outs_0_valid,
      outs_valid(1) => fork10_outs_1_valid,
      outs_ready(0) => fork10_outs_0_ready,
      outs_ready(1) => fork10_outs_1_ready
    );

  mux31 : entity work.mux_dataless(arch) generic map(2, 1)
    port map(
      index => buffer25_outs,
      index_valid => buffer25_outs_valid,
      index_ready => buffer25_outs_ready,
      ins_valid(0) => fork9_outs_1_valid,
      ins_valid(1) => cond_br83_trueOut_valid,
      ins_ready(0) => fork9_outs_1_ready,
      ins_ready(1) => cond_br83_trueOut_ready,
      clk => clk,
      rst => rst,
      outs_valid => mux31_outs_valid,
      outs_ready => mux31_outs_ready
    );

  buffer25 : entity work.tfifo(arch) generic map(5, 1)
    port map(
      ins => fork10_outs_1,
      ins_valid => fork10_outs_1_valid,
      ins_ready => fork10_outs_1_ready,
      clk => clk,
      rst => rst,
      outs => buffer25_outs,
      outs_valid => buffer25_outs_valid,
      outs_ready => buffer25_outs_ready
    );

  buffer32 : entity work.oehb_dataless(arch)
    port map(
      ins_valid => mux31_outs_valid,
      ins_ready => mux31_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer32_outs_valid,
      outs_ready => buffer32_outs_ready
    );

  buffer33 : entity work.tehb_dataless(arch)
    port map(
      ins_valid => buffer32_outs_valid,
      ins_ready => buffer32_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer33_outs_valid,
      outs_ready => buffer33_outs_ready
    );

  fork11 : entity work.fork_dataless(arch) generic map(3)
    port map(
      ins_valid => buffer33_outs_valid,
      ins_ready => buffer33_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid(0) => fork11_outs_0_valid,
      outs_valid(1) => fork11_outs_1_valid,
      outs_valid(2) => fork11_outs_2_valid,
      outs_ready(0) => fork11_outs_0_ready,
      outs_ready(1) => fork11_outs_1_ready,
      outs_ready(2) => fork11_outs_2_ready
    );

  buffer16 : entity work.oehb_dataless(arch)
    port map(
      ins_valid => mux30_outs_valid,
      ins_ready => mux30_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer16_outs_valid,
      outs_ready => buffer16_outs_ready
    );

  buffer17 : entity work.tehb_dataless(arch)
    port map(
      ins_valid => buffer16_outs_valid,
      ins_ready => buffer16_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer17_outs_valid,
      outs_ready => buffer17_outs_ready
    );

  mux34 : entity work.mux_dataless(arch) generic map(2, 1)
    port map(
      index => buffer26_outs,
      index_valid => buffer26_outs_valid,
      index_ready => buffer26_outs_ready,
      ins_valid(0) => buffer17_outs_valid,
      ins_valid(1) => cond_br84_trueOut_valid,
      ins_ready(0) => buffer17_outs_ready,
      ins_ready(1) => cond_br84_trueOut_ready,
      clk => clk,
      rst => rst,
      outs_valid => mux34_outs_valid,
      outs_ready => mux34_outs_ready
    );

  buffer26 : entity work.tfifo(arch) generic map(5, 1)
    port map(
      ins => fork10_outs_0,
      ins_valid => fork10_outs_0_valid,
      ins_ready => fork10_outs_0_ready,
      clk => clk,
      rst => rst,
      outs => buffer26_outs,
      outs_valid => buffer26_outs_valid,
      outs_ready => buffer26_outs_ready
    );

  mux7 : entity work.mux(arch) generic map(2, 5, 1)
    port map(
      index => fork19_outs_2,
      index_valid => fork19_outs_2_valid,
      index_ready => fork19_outs_2_ready,
      ins(0) => extsi32_outs,
      ins(1) => cond_br6_trueOut,
      ins_valid(0) => extsi32_outs_valid,
      ins_valid(1) => cond_br6_trueOut_valid,
      ins_ready(0) => extsi32_outs_ready,
      ins_ready(1) => cond_br6_trueOut_ready,
      clk => clk,
      rst => rst,
      outs => mux7_outs,
      outs_valid => mux7_outs_valid,
      outs_ready => mux7_outs_ready
    );

  buffer40 : entity work.oehb(arch) generic map(5)
    port map(
      ins => mux7_outs,
      ins_valid => mux7_outs_valid,
      ins_ready => mux7_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer40_outs,
      outs_valid => buffer40_outs_valid,
      outs_ready => buffer40_outs_ready
    );

  buffer42 : entity work.tehb(arch) generic map(5)
    port map(
      ins => buffer40_outs,
      ins_valid => buffer40_outs_valid,
      ins_ready => buffer40_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer42_outs,
      outs_valid => buffer42_outs_valid,
      outs_ready => buffer42_outs_ready
    );

  fork12 : entity work.handshake_fork(arch) generic map(3, 5)
    port map(
      ins => buffer42_outs,
      ins_valid => buffer42_outs_valid,
      ins_ready => buffer42_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork12_outs_0,
      outs(1) => fork12_outs_1,
      outs(2) => fork12_outs_2,
      outs_valid(0) => fork12_outs_0_valid,
      outs_valid(1) => fork12_outs_1_valid,
      outs_valid(2) => fork12_outs_2_valid,
      outs_ready(0) => fork12_outs_0_ready,
      outs_ready(1) => fork12_outs_1_ready,
      outs_ready(2) => fork12_outs_2_ready
    );

  extsi37 : entity work.extsi(arch) generic map(5, 7)
    port map(
      ins => buffer28_outs,
      ins_valid => buffer28_outs_valid,
      ins_ready => buffer28_outs_ready,
      clk => clk,
      rst => rst,
      outs => extsi37_outs,
      outs_valid => extsi37_outs_valid,
      outs_ready => extsi37_outs_ready
    );

  buffer28 : entity work.tfifo(arch) generic map(2, 5)
    port map(
      ins => fork12_outs_0,
      ins_valid => fork12_outs_0_valid,
      ins_ready => fork12_outs_0_ready,
      clk => clk,
      rst => rst,
      outs => buffer28_outs,
      outs_valid => buffer28_outs_valid,
      outs_ready => buffer28_outs_ready
    );

  extsi38 : entity work.extsi(arch) generic map(5, 6)
    port map(
      ins => fork12_outs_1,
      ins_valid => fork12_outs_1_valid,
      ins_ready => fork12_outs_1_ready,
      clk => clk,
      rst => rst,
      outs => extsi38_outs,
      outs_valid => extsi38_outs_valid,
      outs_ready => extsi38_outs_ready
    );

  extsi39 : entity work.extsi(arch) generic map(5, 32)
    port map(
      ins => fork12_outs_2,
      ins_valid => fork12_outs_2_valid,
      ins_ready => fork12_outs_2_ready,
      clk => clk,
      rst => rst,
      outs => extsi39_outs,
      outs_valid => extsi39_outs_valid,
      outs_ready => extsi39_outs_ready
    );

  fork13 : entity work.handshake_fork(arch) generic map(2, 32)
    port map(
      ins => extsi39_outs,
      ins_valid => extsi39_outs_valid,
      ins_ready => extsi39_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork13_outs_0,
      outs(1) => fork13_outs_1,
      outs_valid(0) => fork13_outs_0_valid,
      outs_valid(1) => fork13_outs_1_valid,
      outs_ready(0) => fork13_outs_0_ready,
      outs_ready(1) => fork13_outs_1_ready
    );

  mux8 : entity work.mux(arch) generic map(2, 32, 1)
    port map(
      index => fork19_outs_3,
      index_valid => fork19_outs_3_valid,
      index_ready => fork19_outs_3_ready,
      ins(0) => buffer19_outs,
      ins(1) => cond_br7_trueOut,
      ins_valid(0) => buffer19_outs_valid,
      ins_valid(1) => cond_br7_trueOut_valid,
      ins_ready(0) => buffer19_outs_ready,
      ins_ready(1) => cond_br7_trueOut_ready,
      clk => clk,
      rst => rst,
      outs => mux8_outs,
      outs_valid => mux8_outs_valid,
      outs_ready => mux8_outs_ready
    );

  buffer45 : entity work.oehb(arch) generic map(32)
    port map(
      ins => mux8_outs,
      ins_valid => mux8_outs_valid,
      ins_ready => mux8_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer45_outs,
      outs_valid => buffer45_outs_valid,
      outs_ready => buffer45_outs_ready
    );

  buffer47 : entity work.tehb(arch) generic map(32)
    port map(
      ins => buffer45_outs,
      ins_valid => buffer45_outs_valid,
      ins_ready => buffer45_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer47_outs,
      outs_valid => buffer47_outs_valid,
      outs_ready => buffer47_outs_ready
    );

  fork14 : entity work.handshake_fork(arch) generic map(2, 32)
    port map(
      ins => buffer47_outs,
      ins_valid => buffer47_outs_valid,
      ins_ready => buffer47_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork14_outs_0,
      outs(1) => fork14_outs_1,
      outs_valid(0) => fork14_outs_0_valid,
      outs_valid(1) => fork14_outs_1_valid,
      outs_ready(0) => fork14_outs_0_ready,
      outs_ready(1) => fork14_outs_1_ready
    );

  mux9 : entity work.mux(arch) generic map(2, 32, 1)
    port map(
      index => fork19_outs_4,
      index_valid => fork19_outs_4_valid,
      index_ready => fork19_outs_4_ready,
      ins(0) => buffer20_outs,
      ins(1) => cond_br8_trueOut,
      ins_valid(0) => buffer20_outs_valid,
      ins_valid(1) => cond_br8_trueOut_valid,
      ins_ready(0) => buffer20_outs_ready,
      ins_ready(1) => cond_br8_trueOut_ready,
      clk => clk,
      rst => rst,
      outs => mux9_outs,
      outs_valid => mux9_outs_valid,
      outs_ready => mux9_outs_ready
    );

  mux10 : entity work.mux(arch) generic map(2, 5, 1)
    port map(
      index => fork19_outs_0,
      index_valid => fork19_outs_0_valid,
      index_ready => fork19_outs_0_ready,
      ins(0) => fork4_outs_0,
      ins(1) => cond_br9_trueOut,
      ins_valid(0) => fork4_outs_0_valid,
      ins_valid(1) => cond_br9_trueOut_valid,
      ins_ready(0) => fork4_outs_0_ready,
      ins_ready(1) => cond_br9_trueOut_ready,
      clk => clk,
      rst => rst,
      outs => mux10_outs,
      outs_valid => mux10_outs_valid,
      outs_ready => mux10_outs_ready
    );

  buffer72 : entity work.oehb(arch) generic map(5)
    port map(
      ins => mux10_outs,
      ins_valid => mux10_outs_valid,
      ins_ready => mux10_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer72_outs,
      outs_valid => buffer72_outs_valid,
      outs_ready => buffer72_outs_ready
    );

  buffer73 : entity work.tehb(arch) generic map(5)
    port map(
      ins => buffer72_outs,
      ins_valid => buffer72_outs_valid,
      ins_ready => buffer72_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer73_outs,
      outs_valid => buffer73_outs_valid,
      outs_ready => buffer73_outs_ready
    );

  fork15 : entity work.handshake_fork(arch) generic map(2, 5)
    port map(
      ins => buffer73_outs,
      ins_valid => buffer73_outs_valid,
      ins_ready => buffer73_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork15_outs_0,
      outs(1) => fork15_outs_1,
      outs_valid(0) => fork15_outs_0_valid,
      outs_valid(1) => fork15_outs_1_valid,
      outs_ready(0) => fork15_outs_0_ready,
      outs_ready(1) => fork15_outs_1_ready
    );

  extsi40 : entity work.extsi(arch) generic map(5, 32)
    port map(
      ins => buffer34_outs,
      ins_valid => buffer34_outs_valid,
      ins_ready => buffer34_outs_ready,
      clk => clk,
      rst => rst,
      outs => extsi40_outs,
      outs_valid => extsi40_outs_valid,
      outs_ready => extsi40_outs_ready
    );

  buffer34 : entity work.tfifo(arch) generic map(1, 5)
    port map(
      ins => fork15_outs_1,
      ins_valid => fork15_outs_1_valid,
      ins_ready => fork15_outs_1_ready,
      clk => clk,
      rst => rst,
      outs => buffer34_outs,
      outs_valid => buffer34_outs_valid,
      outs_ready => buffer34_outs_ready
    );

  fork16 : entity work.handshake_fork(arch) generic map(6, 32)
    port map(
      ins => extsi40_outs,
      ins_valid => extsi40_outs_valid,
      ins_ready => extsi40_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork16_outs_0,
      outs(1) => fork16_outs_1,
      outs(2) => fork16_outs_2,
      outs(3) => fork16_outs_3,
      outs(4) => fork16_outs_4,
      outs(5) => fork16_outs_5,
      outs_valid(0) => fork16_outs_0_valid,
      outs_valid(1) => fork16_outs_1_valid,
      outs_valid(2) => fork16_outs_2_valid,
      outs_valid(3) => fork16_outs_3_valid,
      outs_valid(4) => fork16_outs_4_valid,
      outs_valid(5) => fork16_outs_5_valid,
      outs_ready(0) => fork16_outs_0_ready,
      outs_ready(1) => fork16_outs_1_ready,
      outs_ready(2) => fork16_outs_2_ready,
      outs_ready(3) => fork16_outs_3_ready,
      outs_ready(4) => fork16_outs_4_ready,
      outs_ready(5) => fork16_outs_5_ready
    );

  mux11 : entity work.mux(arch) generic map(2, 5, 1)
    port map(
      index => buffer35_outs,
      index_valid => buffer35_outs_valid,
      index_ready => buffer35_outs_ready,
      ins(0) => fork3_outs_1,
      ins(1) => cond_br10_trueOut,
      ins_valid(0) => fork3_outs_1_valid,
      ins_valid(1) => cond_br10_trueOut_valid,
      ins_ready(0) => fork3_outs_1_ready,
      ins_ready(1) => cond_br10_trueOut_ready,
      clk => clk,
      rst => rst,
      outs => mux11_outs,
      outs_valid => mux11_outs_valid,
      outs_ready => mux11_outs_ready
    );

  buffer35 : entity work.tfifo(arch) generic map(1, 1)
    port map(
      ins => fork19_outs_1,
      ins_valid => fork19_outs_1_valid,
      ins_ready => fork19_outs_1_ready,
      clk => clk,
      rst => rst,
      outs => buffer35_outs,
      outs_valid => buffer35_outs_valid,
      outs_ready => buffer35_outs_ready
    );

  buffer74 : entity work.oehb(arch) generic map(5)
    port map(
      ins => mux11_outs,
      ins_valid => mux11_outs_valid,
      ins_ready => mux11_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer74_outs,
      outs_valid => buffer74_outs_valid,
      outs_ready => buffer74_outs_ready
    );

  buffer77 : entity work.tehb(arch) generic map(5)
    port map(
      ins => buffer74_outs,
      ins_valid => buffer74_outs_valid,
      ins_ready => buffer74_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer77_outs,
      outs_valid => buffer77_outs_valid,
      outs_ready => buffer77_outs_ready
    );

  fork17 : entity work.handshake_fork(arch) generic map(3, 5)
    port map(
      ins => buffer77_outs,
      ins_valid => buffer77_outs_valid,
      ins_ready => buffer77_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork17_outs_0,
      outs(1) => fork17_outs_1,
      outs(2) => fork17_outs_2,
      outs_valid(0) => fork17_outs_0_valid,
      outs_valid(1) => fork17_outs_1_valid,
      outs_valid(2) => fork17_outs_2_valid,
      outs_ready(0) => fork17_outs_0_ready,
      outs_ready(1) => fork17_outs_1_ready,
      outs_ready(2) => fork17_outs_2_ready
    );

  extsi41 : entity work.extsi(arch) generic map(5, 7)
    port map(
      ins => buffer36_outs,
      ins_valid => buffer36_outs_valid,
      ins_ready => buffer36_outs_ready,
      clk => clk,
      rst => rst,
      outs => extsi41_outs,
      outs_valid => extsi41_outs_valid,
      outs_ready => extsi41_outs_ready
    );

  buffer36 : entity work.tfifo(arch) generic map(1, 5)
    port map(
      ins => fork17_outs_0,
      ins_valid => fork17_outs_0_valid,
      ins_ready => fork17_outs_0_ready,
      clk => clk,
      rst => rst,
      outs => buffer36_outs,
      outs_valid => buffer36_outs_valid,
      outs_ready => buffer36_outs_ready
    );

  extsi42 : entity work.extsi(arch) generic map(5, 32)
    port map(
      ins => fork17_outs_2,
      ins_valid => fork17_outs_2_valid,
      ins_ready => fork17_outs_2_ready,
      clk => clk,
      rst => rst,
      outs => extsi42_outs,
      outs_valid => extsi42_outs_valid,
      outs_ready => extsi42_outs_ready
    );

  fork18 : entity work.handshake_fork(arch) generic map(2, 32)
    port map(
      ins => extsi42_outs,
      ins_valid => extsi42_outs_valid,
      ins_ready => extsi42_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork18_outs_0,
      outs(1) => fork18_outs_1,
      outs_valid(0) => fork18_outs_0_valid,
      outs_valid(1) => fork18_outs_1_valid,
      outs_ready(0) => fork18_outs_0_ready,
      outs_ready(1) => fork18_outs_1_ready
    );

  control_merge2 : entity work.control_merge_dataless(arch) generic map(2, 1)
    port map(
      ins_valid(0) => fork7_outs_2_valid,
      ins_valid(1) => cond_br11_trueOut_valid,
      ins_ready(0) => fork7_outs_2_ready,
      ins_ready(1) => cond_br11_trueOut_ready,
      clk => clk,
      rst => rst,
      outs_valid => control_merge2_outs_valid,
      outs_ready => control_merge2_outs_ready,
      index => control_merge2_index,
      index_valid => control_merge2_index_valid,
      index_ready => control_merge2_index_ready
    );

  fork19 : entity work.handshake_fork(arch) generic map(5, 1)
    port map(
      ins => control_merge2_index,
      ins_valid => control_merge2_index_valid,
      ins_ready => control_merge2_index_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork19_outs_0,
      outs(1) => fork19_outs_1,
      outs(2) => fork19_outs_2,
      outs(3) => fork19_outs_3,
      outs(4) => fork19_outs_4,
      outs_valid(0) => fork19_outs_0_valid,
      outs_valid(1) => fork19_outs_1_valid,
      outs_valid(2) => fork19_outs_2_valid,
      outs_valid(3) => fork19_outs_3_valid,
      outs_valid(4) => fork19_outs_4_valid,
      outs_ready(0) => fork19_outs_0_ready,
      outs_ready(1) => fork19_outs_1_ready,
      outs_ready(2) => fork19_outs_2_ready,
      outs_ready(3) => fork19_outs_3_ready,
      outs_ready(4) => fork19_outs_4_ready
    );

  fork20 : entity work.fork_dataless(arch) generic map(2)
    port map(
      ins_valid => control_merge2_outs_valid,
      ins_ready => control_merge2_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid(0) => fork20_outs_0_valid,
      outs_valid(1) => fork20_outs_1_valid,
      outs_ready(0) => fork20_outs_0_ready,
      outs_ready(1) => fork20_outs_1_ready
    );

  constant35 : entity work.handshake_constant_1(arch) generic map(2)
    port map(
      ctrl_valid => fork20_outs_0_valid,
      ctrl_ready => fork20_outs_0_ready,
      clk => clk,
      rst => rst,
      outs => constant35_outs,
      outs_valid => constant35_outs_valid,
      outs_ready => constant35_outs_ready
    );

  extsi7 : entity work.extsi(arch) generic map(2, 32)
    port map(
      ins => constant35_outs,
      ins_valid => constant35_outs_valid,
      ins_ready => constant35_outs_ready,
      clk => clk,
      rst => rst,
      outs => extsi7_outs,
      outs_valid => extsi7_outs_valid,
      outs_ready => extsi7_outs_ready
    );

  source2 : entity work.source(arch)
    port map(
      clk => clk,
      rst => rst,
      outs_valid => source2_outs_valid,
      outs_ready => source2_outs_ready
    );

  constant36 : entity work.handshake_constant_3(arch) generic map(5)
    port map(
      ctrl_valid => source2_outs_valid,
      ctrl_ready => source2_outs_ready,
      clk => clk,
      rst => rst,
      outs => constant36_outs,
      outs_valid => constant36_outs_valid,
      outs_ready => constant36_outs_ready
    );

  extsi43 : entity work.extsi(arch) generic map(5, 6)
    port map(
      ins => constant36_outs,
      ins_valid => constant36_outs_valid,
      ins_ready => constant36_outs_ready,
      clk => clk,
      rst => rst,
      outs => extsi43_outs,
      outs_valid => extsi43_outs_valid,
      outs_ready => extsi43_outs_ready
    );

  source3 : entity work.source(arch)
    port map(
      clk => clk,
      rst => rst,
      outs_valid => source3_outs_valid,
      outs_ready => source3_outs_ready
    );

  constant37 : entity work.handshake_constant_1(arch) generic map(2)
    port map(
      ctrl_valid => source3_outs_valid,
      ctrl_ready => source3_outs_ready,
      clk => clk,
      rst => rst,
      outs => constant37_outs,
      outs_valid => constant37_outs_valid,
      outs_ready => constant37_outs_ready
    );

  fork21 : entity work.handshake_fork(arch) generic map(2, 2)
    port map(
      ins => constant37_outs,
      ins_valid => constant37_outs_valid,
      ins_ready => constant37_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork21_outs_0,
      outs(1) => fork21_outs_1,
      outs_valid(0) => fork21_outs_0_valid,
      outs_valid(1) => fork21_outs_1_valid,
      outs_ready(0) => fork21_outs_0_ready,
      outs_ready(1) => fork21_outs_1_ready
    );

  extsi44 : entity work.extsi(arch) generic map(2, 6)
    port map(
      ins => buffer38_outs,
      ins_valid => buffer38_outs_valid,
      ins_ready => buffer38_outs_ready,
      clk => clk,
      rst => rst,
      outs => extsi44_outs,
      outs_valid => extsi44_outs_valid,
      outs_ready => extsi44_outs_ready
    );

  buffer38 : entity work.tfifo(arch) generic map(1, 2)
    port map(
      ins => fork21_outs_0,
      ins_valid => fork21_outs_0_valid,
      ins_ready => fork21_outs_0_ready,
      clk => clk,
      rst => rst,
      outs => buffer38_outs,
      outs_valid => buffer38_outs_valid,
      outs_ready => buffer38_outs_ready
    );

  extsi9 : entity work.extsi(arch) generic map(2, 32)
    port map(
      ins => buffer39_outs,
      ins_valid => buffer39_outs_valid,
      ins_ready => buffer39_outs_ready,
      clk => clk,
      rst => rst,
      outs => extsi9_outs,
      outs_valid => extsi9_outs_valid,
      outs_ready => extsi9_outs_ready
    );

  buffer39 : entity work.tfifo(arch) generic map(2, 2)
    port map(
      ins => fork21_outs_1,
      ins_valid => fork21_outs_1_valid,
      ins_ready => fork21_outs_1_ready,
      clk => clk,
      rst => rst,
      outs => buffer39_outs,
      outs_valid => buffer39_outs_valid,
      outs_ready => buffer39_outs_ready
    );

  fork22 : entity work.handshake_fork(arch) generic map(4, 32)
    port map(
      ins => extsi9_outs,
      ins_valid => extsi9_outs_valid,
      ins_ready => extsi9_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork22_outs_0,
      outs(1) => fork22_outs_1,
      outs(2) => fork22_outs_2,
      outs(3) => fork22_outs_3,
      outs_valid(0) => fork22_outs_0_valid,
      outs_valid(1) => fork22_outs_1_valid,
      outs_valid(2) => fork22_outs_2_valid,
      outs_valid(3) => fork22_outs_3_valid,
      outs_ready(0) => fork22_outs_0_ready,
      outs_ready(1) => fork22_outs_1_ready,
      outs_ready(2) => fork22_outs_2_ready,
      outs_ready(3) => fork22_outs_3_ready
    );

  source4 : entity work.source(arch)
    port map(
      clk => clk,
      rst => rst,
      outs_valid => source4_outs_valid,
      outs_ready => source4_outs_ready
    );

  constant38 : entity work.handshake_constant_2(arch) generic map(3)
    port map(
      ctrl_valid => source4_outs_valid,
      ctrl_ready => source4_outs_ready,
      clk => clk,
      rst => rst,
      outs => constant38_outs,
      outs_valid => constant38_outs_valid,
      outs_ready => constant38_outs_ready
    );

  extsi10 : entity work.extsi(arch) generic map(3, 32)
    port map(
      ins => constant38_outs,
      ins_valid => constant38_outs_valid,
      ins_ready => constant38_outs_ready,
      clk => clk,
      rst => rst,
      outs => extsi10_outs,
      outs_valid => extsi10_outs_valid,
      outs_ready => extsi10_outs_ready
    );

  fork23 : entity work.handshake_fork(arch) generic map(4, 32)
    port map(
      ins => extsi10_outs,
      ins_valid => extsi10_outs_valid,
      ins_ready => extsi10_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork23_outs_0,
      outs(1) => fork23_outs_1,
      outs(2) => fork23_outs_2,
      outs(3) => fork23_outs_3,
      outs_valid(0) => fork23_outs_0_valid,
      outs_valid(1) => fork23_outs_1_valid,
      outs_valid(2) => fork23_outs_2_valid,
      outs_valid(3) => fork23_outs_3_valid,
      outs_ready(0) => fork23_outs_0_ready,
      outs_ready(1) => fork23_outs_1_ready,
      outs_ready(2) => fork23_outs_2_ready,
      outs_ready(3) => fork23_outs_3_ready
    );

  shli2 : entity work.shli(arch) generic map(32)
    port map(
      lhs => buffer41_outs,
      lhs_valid => buffer41_outs_valid,
      lhs_ready => buffer41_outs_ready,
      rhs => fork22_outs_0,
      rhs_valid => fork22_outs_0_valid,
      rhs_ready => fork22_outs_0_ready,
      clk => clk,
      rst => rst,
      result => shli2_result,
      result_valid => shli2_result_valid,
      result_ready => shli2_result_ready
    );

  buffer41 : entity work.tfifo(arch) generic map(1, 32)
    port map(
      ins => fork16_outs_0,
      ins_valid => fork16_outs_0_valid,
      ins_ready => fork16_outs_0_ready,
      clk => clk,
      rst => rst,
      outs => buffer41_outs,
      outs_valid => buffer41_outs_valid,
      outs_ready => buffer41_outs_ready
    );

  buffer81 : entity work.oehb(arch) generic map(32)
    port map(
      ins => shli2_result,
      ins_valid => shli2_result_valid,
      ins_ready => shli2_result_ready,
      clk => clk,
      rst => rst,
      outs => buffer81_outs,
      outs_valid => buffer81_outs_valid,
      outs_ready => buffer81_outs_ready
    );

  trunci2 : entity work.trunci(arch) generic map(32, 7)
    port map(
      ins => buffer81_outs,
      ins_valid => buffer81_outs_valid,
      ins_ready => buffer81_outs_ready,
      clk => clk,
      rst => rst,
      outs => trunci2_outs,
      outs_valid => trunci2_outs_valid,
      outs_ready => trunci2_outs_ready
    );

  shli3 : entity work.shli(arch) generic map(32)
    port map(
      lhs => buffer43_outs,
      lhs_valid => buffer43_outs_valid,
      lhs_ready => buffer43_outs_ready,
      rhs => fork23_outs_0,
      rhs_valid => fork23_outs_0_valid,
      rhs_ready => fork23_outs_0_ready,
      clk => clk,
      rst => rst,
      result => shli3_result,
      result_valid => shli3_result_valid,
      result_ready => shli3_result_ready
    );

  buffer43 : entity work.tfifo(arch) generic map(1, 32)
    port map(
      ins => fork16_outs_1,
      ins_valid => fork16_outs_1_valid,
      ins_ready => fork16_outs_1_ready,
      clk => clk,
      rst => rst,
      outs => buffer43_outs,
      outs_valid => buffer43_outs_valid,
      outs_ready => buffer43_outs_ready
    );

  buffer82 : entity work.oehb(arch) generic map(32)
    port map(
      ins => shli3_result,
      ins_valid => shli3_result_valid,
      ins_ready => shli3_result_ready,
      clk => clk,
      rst => rst,
      outs => buffer82_outs,
      outs_valid => buffer82_outs_valid,
      outs_ready => buffer82_outs_ready
    );

  trunci3 : entity work.trunci(arch) generic map(32, 7)
    port map(
      ins => buffer82_outs,
      ins_valid => buffer82_outs_valid,
      ins_ready => buffer82_outs_ready,
      clk => clk,
      rst => rst,
      outs => trunci3_outs,
      outs_valid => trunci3_outs_valid,
      outs_ready => trunci3_outs_ready
    );

  addi20 : entity work.addi(arch) generic map(7)
    port map(
      lhs => trunci2_outs,
      lhs_valid => trunci2_outs_valid,
      lhs_ready => trunci2_outs_ready,
      rhs => trunci3_outs,
      rhs_valid => trunci3_outs_valid,
      rhs_ready => trunci3_outs_ready,
      clk => clk,
      rst => rst,
      result => addi20_result,
      result_valid => addi20_result_valid,
      result_ready => addi20_result_ready
    );

  buffer83 : entity work.oehb(arch) generic map(7)
    port map(
      ins => addi20_result,
      ins_valid => addi20_result_valid,
      ins_ready => addi20_result_ready,
      clk => clk,
      rst => rst,
      outs => buffer83_outs,
      outs_valid => buffer83_outs_valid,
      outs_ready => buffer83_outs_ready
    );

  addi3 : entity work.addi(arch) generic map(7)
    port map(
      lhs => extsi37_outs,
      lhs_valid => extsi37_outs_valid,
      lhs_ready => extsi37_outs_ready,
      rhs => buffer83_outs,
      rhs_valid => buffer83_outs_valid,
      rhs_ready => buffer83_outs_ready,
      clk => clk,
      rst => rst,
      result => addi3_result,
      result_valid => addi3_result_valid,
      result_ready => addi3_result_ready
    );

  load0 : entity work.load(arch) generic map(32, 7)
    port map(
      addrIn => addi3_result,
      addrIn_valid => addi3_result_valid,
      addrIn_ready => addi3_result_ready,
      dataFromMem => mem_controller6_ldData_0,
      dataFromMem_valid => mem_controller6_ldData_0_valid,
      dataFromMem_ready => mem_controller6_ldData_0_ready,
      clk => clk,
      rst => rst,
      addrOut => load0_addrOut,
      addrOut_valid => load0_addrOut_valid,
      addrOut_ready => load0_addrOut_ready,
      dataOut => load0_dataOut,
      dataOut_valid => load0_dataOut_valid,
      dataOut_ready => load0_dataOut_ready
    );

  muli0 : entity work.muli(arch) generic map(32)
    port map(
      lhs => buffer44_outs,
      lhs_valid => buffer44_outs_valid,
      lhs_ready => buffer44_outs_ready,
      rhs => load0_dataOut,
      rhs_valid => load0_dataOut_valid,
      rhs_ready => load0_dataOut_ready,
      clk => clk,
      rst => rst,
      result => muli0_result,
      result_valid => muli0_result_valid,
      result_ready => muli0_result_ready
    );

  buffer44 : entity work.tfifo(arch) generic map(1, 32)
    port map(
      ins => fork14_outs_1,
      ins_valid => fork14_outs_1_valid,
      ins_ready => fork14_outs_1_ready,
      clk => clk,
      rst => rst,
      outs => buffer44_outs,
      outs_valid => buffer44_outs_valid,
      outs_ready => buffer44_outs_ready
    );

  shli4 : entity work.shli(arch) generic map(32)
    port map(
      lhs => buffer46_outs,
      lhs_valid => buffer46_outs_valid,
      lhs_ready => buffer46_outs_ready,
      rhs => fork22_outs_1,
      rhs_valid => fork22_outs_1_valid,
      rhs_ready => fork22_outs_1_ready,
      clk => clk,
      rst => rst,
      result => shli4_result,
      result_valid => shli4_result_valid,
      result_ready => shli4_result_ready
    );

  buffer46 : entity work.tfifo(arch) generic map(2, 32)
    port map(
      ins => fork13_outs_0,
      ins_valid => fork13_outs_0_valid,
      ins_ready => fork13_outs_0_ready,
      clk => clk,
      rst => rst,
      outs => buffer46_outs,
      outs_valid => buffer46_outs_valid,
      outs_ready => buffer46_outs_ready
    );

  buffer84 : entity work.oehb(arch) generic map(32)
    port map(
      ins => shli4_result,
      ins_valid => shli4_result_valid,
      ins_ready => shli4_result_ready,
      clk => clk,
      rst => rst,
      outs => buffer84_outs,
      outs_valid => buffer84_outs_valid,
      outs_ready => buffer84_outs_ready
    );

  trunci4 : entity work.trunci(arch) generic map(32, 7)
    port map(
      ins => buffer84_outs,
      ins_valid => buffer84_outs_valid,
      ins_ready => buffer84_outs_ready,
      clk => clk,
      rst => rst,
      outs => trunci4_outs,
      outs_valid => trunci4_outs_valid,
      outs_ready => trunci4_outs_ready
    );

  shli5 : entity work.shli(arch) generic map(32)
    port map(
      lhs => buffer48_outs,
      lhs_valid => buffer48_outs_valid,
      lhs_ready => buffer48_outs_ready,
      rhs => fork23_outs_1,
      rhs_valid => fork23_outs_1_valid,
      rhs_ready => fork23_outs_1_ready,
      clk => clk,
      rst => rst,
      result => shli5_result,
      result_valid => shli5_result_valid,
      result_ready => shli5_result_ready
    );

  buffer48 : entity work.tfifo(arch) generic map(2, 32)
    port map(
      ins => fork13_outs_1,
      ins_valid => fork13_outs_1_valid,
      ins_ready => fork13_outs_1_ready,
      clk => clk,
      rst => rst,
      outs => buffer48_outs,
      outs_valid => buffer48_outs_valid,
      outs_ready => buffer48_outs_ready
    );

  buffer85 : entity work.oehb(arch) generic map(32)
    port map(
      ins => shli5_result,
      ins_valid => shli5_result_valid,
      ins_ready => shli5_result_ready,
      clk => clk,
      rst => rst,
      outs => buffer85_outs,
      outs_valid => buffer85_outs_valid,
      outs_ready => buffer85_outs_ready
    );

  trunci5 : entity work.trunci(arch) generic map(32, 7)
    port map(
      ins => buffer85_outs,
      ins_valid => buffer85_outs_valid,
      ins_ready => buffer85_outs_ready,
      clk => clk,
      rst => rst,
      outs => trunci5_outs,
      outs_valid => trunci5_outs_valid,
      outs_ready => trunci5_outs_ready
    );

  addi21 : entity work.addi(arch) generic map(7)
    port map(
      lhs => trunci4_outs,
      lhs_valid => trunci4_outs_valid,
      lhs_ready => trunci4_outs_ready,
      rhs => trunci5_outs,
      rhs_valid => trunci5_outs_valid,
      rhs_ready => trunci5_outs_ready,
      clk => clk,
      rst => rst,
      result => addi21_result,
      result_valid => addi21_result_valid,
      result_ready => addi21_result_ready
    );

  buffer86 : entity work.oehb(arch) generic map(7)
    port map(
      ins => addi21_result,
      ins_valid => addi21_result_valid,
      ins_ready => addi21_result_ready,
      clk => clk,
      rst => rst,
      outs => buffer86_outs,
      outs_valid => buffer86_outs_valid,
      outs_ready => buffer86_outs_ready
    );

  addi4 : entity work.addi(arch) generic map(7)
    port map(
      lhs => extsi41_outs,
      lhs_valid => extsi41_outs_valid,
      lhs_ready => extsi41_outs_ready,
      rhs => buffer86_outs,
      rhs_valid => buffer86_outs_valid,
      rhs_ready => buffer86_outs_ready,
      clk => clk,
      rst => rst,
      result => addi4_result,
      result_valid => addi4_result_valid,
      result_ready => addi4_result_ready
    );

  load1 : entity work.load(arch) generic map(32, 7)
    port map(
      addrIn => addi4_result,
      addrIn_valid => addi4_result_valid,
      addrIn_ready => addi4_result_ready,
      dataFromMem => mem_controller5_ldData_0,
      dataFromMem_valid => mem_controller5_ldData_0_valid,
      dataFromMem_ready => mem_controller5_ldData_0_ready,
      clk => clk,
      rst => rst,
      addrOut => load1_addrOut,
      addrOut_valid => load1_addrOut_valid,
      addrOut_ready => load1_addrOut_ready,
      dataOut => load1_dataOut,
      dataOut_valid => load1_dataOut_valid,
      dataOut_ready => load1_dataOut_ready
    );

  muli1 : entity work.muli(arch) generic map(32)
    port map(
      lhs => muli0_result,
      lhs_valid => muli0_result_valid,
      lhs_ready => muli0_result_ready,
      rhs => load1_dataOut,
      rhs_valid => load1_dataOut_valid,
      rhs_ready => load1_dataOut_ready,
      clk => clk,
      rst => rst,
      result => muli1_result,
      result_valid => muli1_result_valid,
      result_ready => muli1_result_ready
    );

  shli6 : entity work.shli(arch) generic map(32)
    port map(
      lhs => buffer50_outs,
      lhs_valid => buffer50_outs_valid,
      lhs_ready => buffer50_outs_ready,
      rhs => buffer49_outs,
      rhs_valid => buffer49_outs_valid,
      rhs_ready => buffer49_outs_ready,
      clk => clk,
      rst => rst,
      result => shli6_result,
      result_valid => shli6_result_valid,
      result_ready => shli6_result_ready
    );

  buffer49 : entity work.tfifo(arch) generic map(5, 32)
    port map(
      ins => fork22_outs_2,
      ins_valid => fork22_outs_2_valid,
      ins_ready => fork22_outs_2_ready,
      clk => clk,
      rst => rst,
      outs => buffer49_outs,
      outs_valid => buffer49_outs_valid,
      outs_ready => buffer49_outs_ready
    );

  buffer50 : entity work.tfifo(arch) generic map(5, 32)
    port map(
      ins => fork16_outs_2,
      ins_valid => fork16_outs_2_valid,
      ins_ready => fork16_outs_2_ready,
      clk => clk,
      rst => rst,
      outs => buffer50_outs,
      outs_valid => buffer50_outs_valid,
      outs_ready => buffer50_outs_ready
    );

  shli7 : entity work.shli(arch) generic map(32)
    port map(
      lhs => buffer52_outs,
      lhs_valid => buffer52_outs_valid,
      lhs_ready => buffer52_outs_ready,
      rhs => buffer51_outs,
      rhs_valid => buffer51_outs_valid,
      rhs_ready => buffer51_outs_ready,
      clk => clk,
      rst => rst,
      result => shli7_result,
      result_valid => shli7_result_valid,
      result_ready => shli7_result_ready
    );

  buffer51 : entity work.tfifo(arch) generic map(5, 32)
    port map(
      ins => fork23_outs_2,
      ins_valid => fork23_outs_2_valid,
      ins_ready => fork23_outs_2_ready,
      clk => clk,
      rst => rst,
      outs => buffer51_outs,
      outs_valid => buffer51_outs_valid,
      outs_ready => buffer51_outs_ready
    );

  buffer52 : entity work.tfifo(arch) generic map(5, 32)
    port map(
      ins => fork16_outs_3,
      ins_valid => fork16_outs_3_valid,
      ins_ready => fork16_outs_3_ready,
      clk => clk,
      rst => rst,
      outs => buffer52_outs,
      outs_valid => buffer52_outs_valid,
      outs_ready => buffer52_outs_ready
    );

  buffer87 : entity work.oehb(arch) generic map(32)
    port map(
      ins => shli6_result,
      ins_valid => shli6_result_valid,
      ins_ready => shli6_result_ready,
      clk => clk,
      rst => rst,
      outs => buffer87_outs,
      outs_valid => buffer87_outs_valid,
      outs_ready => buffer87_outs_ready
    );

  buffer88 : entity work.oehb(arch) generic map(32)
    port map(
      ins => shli7_result,
      ins_valid => shli7_result_valid,
      ins_ready => shli7_result_ready,
      clk => clk,
      rst => rst,
      outs => buffer88_outs,
      outs_valid => buffer88_outs_valid,
      outs_ready => buffer88_outs_ready
    );

  addi22 : entity work.addi(arch) generic map(32)
    port map(
      lhs => buffer87_outs,
      lhs_valid => buffer87_outs_valid,
      lhs_ready => buffer87_outs_ready,
      rhs => buffer88_outs,
      rhs_valid => buffer88_outs_valid,
      rhs_ready => buffer88_outs_ready,
      clk => clk,
      rst => rst,
      result => addi22_result,
      result_valid => addi22_result_valid,
      result_ready => addi22_result_ready
    );

  buffer92 : entity work.oehb(arch) generic map(32)
    port map(
      ins => addi22_result,
      ins_valid => addi22_result_valid,
      ins_ready => addi22_result_ready,
      clk => clk,
      rst => rst,
      outs => buffer92_outs,
      outs_valid => buffer92_outs_valid,
      outs_ready => buffer92_outs_ready
    );

  addi5 : entity work.addi(arch) generic map(32)
    port map(
      lhs => buffer53_outs,
      lhs_valid => buffer53_outs_valid,
      lhs_ready => buffer53_outs_ready,
      rhs => buffer92_outs,
      rhs_valid => buffer92_outs_valid,
      rhs_ready => buffer92_outs_ready,
      clk => clk,
      rst => rst,
      result => addi5_result,
      result_valid => addi5_result_valid,
      result_ready => addi5_result_ready
    );

  buffer53 : entity work.tfifo(arch) generic map(4, 32)
    port map(
      ins => fork18_outs_0,
      ins_valid => fork18_outs_0_valid,
      ins_ready => fork18_outs_0_ready,
      clk => clk,
      rst => rst,
      outs => buffer53_outs,
      outs_valid => buffer53_outs_valid,
      outs_ready => buffer53_outs_ready
    );

  buffer37 : entity work.tehb_dataless(arch)
    port map(
      ins_valid => mux34_outs_valid,
      ins_ready => mux34_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer37_outs_valid,
      outs_ready => buffer37_outs_ready
    );

  gate0 : entity work.gate(arch) generic map(3, 32)
    port map(
      ins(0) => addi5_result,
      ins_valid(0) => addi5_result_valid,
      ins_valid(1) => fork11_outs_1_valid,
      ins_valid(2) => buffer37_outs_valid,
      ins_ready(0) => addi5_result_ready,
      ins_ready(1) => fork11_outs_1_ready,
      ins_ready(2) => buffer37_outs_ready,
      clk => clk,
      rst => rst,
      outs => gate0_outs,
      outs_valid => gate0_outs_valid,
      outs_ready => gate0_outs_ready
    );

  trunci6 : entity work.trunci(arch) generic map(32, 7)
    port map(
      ins => gate0_outs,
      ins_valid => gate0_outs_valid,
      ins_ready => gate0_outs_ready,
      clk => clk,
      rst => rst,
      outs => trunci6_outs,
      outs_valid => trunci6_outs_valid,
      outs_ready => trunci6_outs_ready
    );

  load2 : entity work.load(arch) generic map(32, 7)
    port map(
      addrIn => trunci6_outs,
      addrIn_valid => trunci6_outs_valid,
      addrIn_ready => trunci6_outs_ready,
      dataFromMem => mem_controller7_ldData_0,
      dataFromMem_valid => mem_controller7_ldData_0_valid,
      dataFromMem_ready => mem_controller7_ldData_0_ready,
      clk => clk,
      rst => rst,
      addrOut => load2_addrOut,
      addrOut_valid => load2_addrOut_valid,
      addrOut_ready => load2_addrOut_ready,
      dataOut => load2_dataOut,
      dataOut_valid => load2_dataOut_valid,
      dataOut_ready => load2_dataOut_ready
    );

  addi0 : entity work.addi(arch) generic map(32)
    port map(
      lhs => load2_dataOut,
      lhs_valid => load2_dataOut_valid,
      lhs_ready => load2_dataOut_ready,
      rhs => muli1_result,
      rhs_valid => muli1_result_valid,
      rhs_ready => muli1_result_ready,
      clk => clk,
      rst => rst,
      result => addi0_result,
      result_valid => addi0_result_valid,
      result_ready => addi0_result_ready
    );

  shli8 : entity work.shli(arch) generic map(32)
    port map(
      lhs => buffer55_outs,
      lhs_valid => buffer55_outs_valid,
      lhs_ready => buffer55_outs_ready,
      rhs => buffer54_outs,
      rhs_valid => buffer54_outs_valid,
      rhs_ready => buffer54_outs_ready,
      clk => clk,
      rst => rst,
      result => shli8_result,
      result_valid => shli8_result_valid,
      result_ready => shli8_result_ready
    );

  buffer54 : entity work.tfifo(arch) generic map(4, 32)
    port map(
      ins => fork22_outs_3,
      ins_valid => fork22_outs_3_valid,
      ins_ready => fork22_outs_3_ready,
      clk => clk,
      rst => rst,
      outs => buffer54_outs,
      outs_valid => buffer54_outs_valid,
      outs_ready => buffer54_outs_ready
    );

  buffer55 : entity work.tfifo(arch) generic map(4, 32)
    port map(
      ins => fork16_outs_4,
      ins_valid => fork16_outs_4_valid,
      ins_ready => fork16_outs_4_ready,
      clk => clk,
      rst => rst,
      outs => buffer55_outs,
      outs_valid => buffer55_outs_valid,
      outs_ready => buffer55_outs_ready
    );

  shli9 : entity work.shli(arch) generic map(32)
    port map(
      lhs => buffer57_outs,
      lhs_valid => buffer57_outs_valid,
      lhs_ready => buffer57_outs_ready,
      rhs => buffer56_outs,
      rhs_valid => buffer56_outs_valid,
      rhs_ready => buffer56_outs_ready,
      clk => clk,
      rst => rst,
      result => shli9_result,
      result_valid => shli9_result_valid,
      result_ready => shli9_result_ready
    );

  buffer56 : entity work.tfifo(arch) generic map(4, 32)
    port map(
      ins => fork23_outs_3,
      ins_valid => fork23_outs_3_valid,
      ins_ready => fork23_outs_3_ready,
      clk => clk,
      rst => rst,
      outs => buffer56_outs,
      outs_valid => buffer56_outs_valid,
      outs_ready => buffer56_outs_ready
    );

  buffer57 : entity work.tfifo(arch) generic map(4, 32)
    port map(
      ins => fork16_outs_5,
      ins_valid => fork16_outs_5_valid,
      ins_ready => fork16_outs_5_ready,
      clk => clk,
      rst => rst,
      outs => buffer57_outs,
      outs_valid => buffer57_outs_valid,
      outs_ready => buffer57_outs_ready
    );

  buffer93 : entity work.oehb(arch) generic map(32)
    port map(
      ins => shli8_result,
      ins_valid => shli8_result_valid,
      ins_ready => shli8_result_ready,
      clk => clk,
      rst => rst,
      outs => buffer93_outs,
      outs_valid => buffer93_outs_valid,
      outs_ready => buffer93_outs_ready
    );

  buffer94 : entity work.oehb(arch) generic map(32)
    port map(
      ins => shli9_result,
      ins_valid => shli9_result_valid,
      ins_ready => shli9_result_ready,
      clk => clk,
      rst => rst,
      outs => buffer94_outs,
      outs_valid => buffer94_outs_valid,
      outs_ready => buffer94_outs_ready
    );

  addi23 : entity work.addi(arch) generic map(32)
    port map(
      lhs => buffer93_outs,
      lhs_valid => buffer93_outs_valid,
      lhs_ready => buffer93_outs_ready,
      rhs => buffer94_outs,
      rhs_valid => buffer94_outs_valid,
      rhs_ready => buffer94_outs_ready,
      clk => clk,
      rst => rst,
      result => addi23_result,
      result_valid => addi23_result_valid,
      result_ready => addi23_result_ready
    );

  buffer99 : entity work.oehb(arch) generic map(32)
    port map(
      ins => addi23_result,
      ins_valid => addi23_result_valid,
      ins_ready => addi23_result_ready,
      clk => clk,
      rst => rst,
      outs => buffer99_outs,
      outs_valid => buffer99_outs_valid,
      outs_ready => buffer99_outs_ready
    );

  addi6 : entity work.addi(arch) generic map(32)
    port map(
      lhs => buffer58_outs,
      lhs_valid => buffer58_outs_valid,
      lhs_ready => buffer58_outs_ready,
      rhs => buffer99_outs,
      rhs_valid => buffer99_outs_valid,
      rhs_ready => buffer99_outs_ready,
      clk => clk,
      rst => rst,
      result => addi6_result,
      result_valid => addi6_result_valid,
      result_ready => addi6_result_ready
    );

  buffer58 : entity work.tfifo(arch) generic map(5, 32)
    port map(
      ins => fork18_outs_1,
      ins_valid => fork18_outs_1_valid,
      ins_ready => fork18_outs_1_ready,
      clk => clk,
      rst => rst,
      outs => buffer58_outs,
      outs_valid => buffer58_outs_valid,
      outs_ready => buffer58_outs_ready
    );

  buffer1 : entity work.tfifo_dataless(arch) generic map(1)
    port map(
      ins_valid => store1_doneOut_valid,
      ins_ready => store1_doneOut_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer1_outs_valid,
      outs_ready => buffer1_outs_ready
    );

  gate1 : entity work.gate(arch) generic map(2, 32)
    port map(
      ins(0) => addi6_result,
      ins_valid(0) => addi6_result_valid,
      ins_valid(1) => fork11_outs_0_valid,
      ins_ready(0) => addi6_result_ready,
      ins_ready(1) => fork11_outs_0_ready,
      clk => clk,
      rst => rst,
      outs => gate1_outs,
      outs_valid => gate1_outs_valid,
      outs_ready => gate1_outs_ready
    );

  trunci7 : entity work.trunci(arch) generic map(32, 7)
    port map(
      ins => gate1_outs,
      ins_valid => gate1_outs_valid,
      ins_ready => gate1_outs_ready,
      clk => clk,
      rst => rst,
      outs => trunci7_outs,
      outs_valid => trunci7_outs_valid,
      outs_ready => trunci7_outs_ready
    );

  store1 : entity work.store(arch) generic map(32, 7)
    port map(
      addrIn => trunci7_outs,
      addrIn_valid => trunci7_outs_valid,
      addrIn_ready => trunci7_outs_ready,
      dataIn => addi0_result,
      dataIn_valid => addi0_result_valid,
      dataIn_ready => addi0_result_ready,
      doneFromMem_valid => mem_controller7_stDone_1_valid,
      doneFromMem_ready => mem_controller7_stDone_1_ready,
      clk => clk,
      rst => rst,
      addrOut => store1_addrOut,
      addrOut_valid => store1_addrOut_valid,
      addrOut_ready => store1_addrOut_ready,
      dataToMem => store1_dataToMem,
      dataToMem_valid => store1_dataToMem_valid,
      dataToMem_ready => store1_dataToMem_ready,
      doneOut_valid => store1_doneOut_valid,
      doneOut_ready => store1_doneOut_ready
    );

  addi13 : entity work.addi(arch) generic map(6)
    port map(
      lhs => extsi38_outs,
      lhs_valid => extsi38_outs_valid,
      lhs_ready => extsi38_outs_ready,
      rhs => extsi44_outs,
      rhs_valid => extsi44_outs_valid,
      rhs_ready => extsi44_outs_ready,
      clk => clk,
      rst => rst,
      result => addi13_result,
      result_valid => addi13_result_valid,
      result_ready => addi13_result_ready
    );

  fork24 : entity work.handshake_fork(arch) generic map(2, 6)
    port map(
      ins => addi13_result,
      ins_valid => addi13_result_valid,
      ins_ready => addi13_result_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork24_outs_0,
      outs(1) => fork24_outs_1,
      outs_valid(0) => fork24_outs_0_valid,
      outs_valid(1) => fork24_outs_1_valid,
      outs_ready(0) => fork24_outs_0_ready,
      outs_ready(1) => fork24_outs_1_ready
    );

  trunci8 : entity work.trunci(arch) generic map(6, 5)
    port map(
      ins => buffer59_outs,
      ins_valid => buffer59_outs_valid,
      ins_ready => buffer59_outs_ready,
      clk => clk,
      rst => rst,
      outs => trunci8_outs,
      outs_valid => trunci8_outs_valid,
      outs_ready => trunci8_outs_ready
    );

  buffer59 : entity work.tfifo(arch) generic map(1, 6)
    port map(
      ins => fork24_outs_0,
      ins_valid => fork24_outs_0_valid,
      ins_ready => fork24_outs_0_ready,
      clk => clk,
      rst => rst,
      outs => buffer59_outs,
      outs_valid => buffer59_outs_valid,
      outs_ready => buffer59_outs_ready
    );

  buffer103 : entity work.oehb(arch) generic map(6)
    port map(
      ins => buffer60_outs,
      ins_valid => buffer60_outs_valid,
      ins_ready => buffer60_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer103_outs,
      outs_valid => buffer103_outs_valid,
      outs_ready => buffer103_outs_ready
    );

  cmpi0 : entity work.handshake_cmpi_0(arch) generic map(6)
    port map(
      lhs => buffer103_outs,
      lhs_valid => buffer103_outs_valid,
      lhs_ready => buffer103_outs_ready,
      rhs => extsi43_outs,
      rhs_valid => extsi43_outs_valid,
      rhs_ready => extsi43_outs_ready,
      clk => clk,
      rst => rst,
      result => cmpi0_result,
      result_valid => cmpi0_result_valid,
      result_ready => cmpi0_result_ready
    );

  buffer60 : entity work.tfifo(arch) generic map(1, 6)
    port map(
      ins => fork24_outs_1,
      ins_valid => fork24_outs_1_valid,
      ins_ready => fork24_outs_1_ready,
      clk => clk,
      rst => rst,
      outs => buffer60_outs,
      outs_valid => buffer60_outs_valid,
      outs_ready => buffer60_outs_ready
    );

  buffer102 : entity work.oehb(arch) generic map(1)
    port map(
      ins => cmpi0_result,
      ins_valid => cmpi0_result_valid,
      ins_ready => cmpi0_result_ready,
      clk => clk,
      rst => rst,
      outs => buffer102_outs,
      outs_valid => buffer102_outs_valid,
      outs_ready => buffer102_outs_ready
    );

  fork25 : entity work.handshake_fork(arch) generic map(9, 1)
    port map(
      ins => buffer102_outs,
      ins_valid => buffer102_outs_valid,
      ins_ready => buffer102_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork25_outs_0,
      outs(1) => fork25_outs_1,
      outs(2) => fork25_outs_2,
      outs(3) => fork25_outs_3,
      outs(4) => fork25_outs_4,
      outs(5) => fork25_outs_5,
      outs(6) => fork25_outs_6,
      outs(7) => fork25_outs_7,
      outs(8) => fork25_outs_8,
      outs_valid(0) => fork25_outs_0_valid,
      outs_valid(1) => fork25_outs_1_valid,
      outs_valid(2) => fork25_outs_2_valid,
      outs_valid(3) => fork25_outs_3_valid,
      outs_valid(4) => fork25_outs_4_valid,
      outs_valid(5) => fork25_outs_5_valid,
      outs_valid(6) => fork25_outs_6_valid,
      outs_valid(7) => fork25_outs_7_valid,
      outs_valid(8) => fork25_outs_8_valid,
      outs_ready(0) => fork25_outs_0_ready,
      outs_ready(1) => fork25_outs_1_ready,
      outs_ready(2) => fork25_outs_2_ready,
      outs_ready(3) => fork25_outs_3_ready,
      outs_ready(4) => fork25_outs_4_ready,
      outs_ready(5) => fork25_outs_5_ready,
      outs_ready(6) => fork25_outs_6_ready,
      outs_ready(7) => fork25_outs_7_ready,
      outs_ready(8) => fork25_outs_8_ready
    );

  cond_br6 : entity work.cond_br(arch) generic map(5)
    port map(
      condition => fork25_outs_0,
      condition_valid => fork25_outs_0_valid,
      condition_ready => fork25_outs_0_ready,
      data => trunci8_outs,
      data_valid => trunci8_outs_valid,
      data_ready => trunci8_outs_ready,
      clk => clk,
      rst => rst,
      trueOut => cond_br6_trueOut,
      trueOut_valid => cond_br6_trueOut_valid,
      trueOut_ready => cond_br6_trueOut_ready,
      falseOut => cond_br6_falseOut,
      falseOut_valid => cond_br6_falseOut_valid,
      falseOut_ready => cond_br6_falseOut_ready
    );

  sink1 : entity work.sink(arch) generic map(5)
    port map(
      ins => cond_br6_falseOut,
      ins_valid => cond_br6_falseOut_valid,
      ins_ready => cond_br6_falseOut_ready,
      clk => clk,
      rst => rst
    );

  cond_br7 : entity work.cond_br(arch) generic map(32)
    port map(
      condition => buffer62_outs,
      condition_valid => buffer62_outs_valid,
      condition_ready => buffer62_outs_ready,
      data => buffer63_outs,
      data_valid => buffer63_outs_valid,
      data_ready => buffer63_outs_ready,
      clk => clk,
      rst => rst,
      trueOut => cond_br7_trueOut,
      trueOut_valid => cond_br7_trueOut_valid,
      trueOut_ready => cond_br7_trueOut_ready,
      falseOut => cond_br7_falseOut,
      falseOut_valid => cond_br7_falseOut_valid,
      falseOut_ready => cond_br7_falseOut_ready
    );

  buffer62 : entity work.tfifo(arch) generic map(1, 1)
    port map(
      ins => fork25_outs_6,
      ins_valid => fork25_outs_6_valid,
      ins_ready => fork25_outs_6_ready,
      clk => clk,
      rst => rst,
      outs => buffer62_outs,
      outs_valid => buffer62_outs_valid,
      outs_ready => buffer62_outs_ready
    );

  buffer63 : entity work.tfifo(arch) generic map(1, 32)
    port map(
      ins => fork14_outs_0,
      ins_valid => fork14_outs_0_valid,
      ins_ready => fork14_outs_0_ready,
      clk => clk,
      rst => rst,
      outs => buffer63_outs,
      outs_valid => buffer63_outs_valid,
      outs_ready => buffer63_outs_ready
    );

  buffer61 : entity work.oehb(arch) generic map(32)
    port map(
      ins => mux9_outs,
      ins_valid => mux9_outs_valid,
      ins_ready => mux9_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer61_outs,
      outs_valid => buffer61_outs_valid,
      outs_ready => buffer61_outs_ready
    );

  buffer67 : entity work.tehb(arch) generic map(32)
    port map(
      ins => buffer61_outs,
      ins_valid => buffer61_outs_valid,
      ins_ready => buffer61_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer67_outs,
      outs_valid => buffer67_outs_valid,
      outs_ready => buffer67_outs_ready
    );

  cond_br8 : entity work.cond_br(arch) generic map(32)
    port map(
      condition => buffer64_outs,
      condition_valid => buffer64_outs_valid,
      condition_ready => buffer64_outs_ready,
      data => buffer67_outs,
      data_valid => buffer67_outs_valid,
      data_ready => buffer67_outs_ready,
      clk => clk,
      rst => rst,
      trueOut => cond_br8_trueOut,
      trueOut_valid => cond_br8_trueOut_valid,
      trueOut_ready => cond_br8_trueOut_ready,
      falseOut => cond_br8_falseOut,
      falseOut_valid => cond_br8_falseOut_valid,
      falseOut_ready => cond_br8_falseOut_ready
    );

  buffer64 : entity work.tfifo(arch) generic map(1, 1)
    port map(
      ins => fork25_outs_7,
      ins_valid => fork25_outs_7_valid,
      ins_ready => fork25_outs_7_ready,
      clk => clk,
      rst => rst,
      outs => buffer64_outs,
      outs_valid => buffer64_outs_valid,
      outs_ready => buffer64_outs_ready
    );

  cond_br9 : entity work.cond_br(arch) generic map(5)
    port map(
      condition => buffer65_outs,
      condition_valid => buffer65_outs_valid,
      condition_ready => buffer65_outs_ready,
      data => buffer66_outs,
      data_valid => buffer66_outs_valid,
      data_ready => buffer66_outs_ready,
      clk => clk,
      rst => rst,
      trueOut => cond_br9_trueOut,
      trueOut_valid => cond_br9_trueOut_valid,
      trueOut_ready => cond_br9_trueOut_ready,
      falseOut => cond_br9_falseOut,
      falseOut_valid => cond_br9_falseOut_valid,
      falseOut_ready => cond_br9_falseOut_ready
    );

  buffer65 : entity work.tfifo(arch) generic map(1, 1)
    port map(
      ins => fork25_outs_1,
      ins_valid => fork25_outs_1_valid,
      ins_ready => fork25_outs_1_ready,
      clk => clk,
      rst => rst,
      outs => buffer65_outs,
      outs_valid => buffer65_outs_valid,
      outs_ready => buffer65_outs_ready
    );

  buffer66 : entity work.tfifo(arch) generic map(1, 5)
    port map(
      ins => fork15_outs_0,
      ins_valid => fork15_outs_0_valid,
      ins_ready => fork15_outs_0_ready,
      clk => clk,
      rst => rst,
      outs => buffer66_outs,
      outs_valid => buffer66_outs_valid,
      outs_ready => buffer66_outs_ready
    );

  cond_br10 : entity work.cond_br(arch) generic map(5)
    port map(
      condition => fork25_outs_2,
      condition_valid => fork25_outs_2_valid,
      condition_ready => fork25_outs_2_ready,
      data => buffer68_outs,
      data_valid => buffer68_outs_valid,
      data_ready => buffer68_outs_ready,
      clk => clk,
      rst => rst,
      trueOut => cond_br10_trueOut,
      trueOut_valid => cond_br10_trueOut_valid,
      trueOut_ready => cond_br10_trueOut_ready,
      falseOut => cond_br10_falseOut,
      falseOut_valid => cond_br10_falseOut_valid,
      falseOut_ready => cond_br10_falseOut_ready
    );

  buffer68 : entity work.tfifo(arch) generic map(1, 5)
    port map(
      ins => fork17_outs_1,
      ins_valid => fork17_outs_1_valid,
      ins_ready => fork17_outs_1_ready,
      clk => clk,
      rst => rst,
      outs => buffer68_outs,
      outs_valid => buffer68_outs_valid,
      outs_ready => buffer68_outs_ready
    );

  buffer79 : entity work.oehb_dataless(arch)
    port map(
      ins_valid => fork20_outs_1_valid,
      ins_ready => fork20_outs_1_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer79_outs_valid,
      outs_ready => buffer79_outs_ready
    );

  cond_br11 : entity work.cond_br_dataless(arch)
    port map(
      condition => buffer69_outs,
      condition_valid => buffer69_outs_valid,
      condition_ready => buffer69_outs_ready,
      data_valid => buffer79_outs_valid,
      data_ready => buffer79_outs_ready,
      clk => clk,
      rst => rst,
      trueOut_valid => cond_br11_trueOut_valid,
      trueOut_ready => cond_br11_trueOut_ready,
      falseOut_valid => cond_br11_falseOut_valid,
      falseOut_ready => cond_br11_falseOut_ready
    );

  buffer69 : entity work.tfifo(arch) generic map(1, 1)
    port map(
      ins => fork25_outs_8,
      ins_valid => fork25_outs_8_valid,
      ins_ready => fork25_outs_8_ready,
      clk => clk,
      rst => rst,
      outs => buffer69_outs,
      outs_valid => buffer69_outs_valid,
      outs_ready => buffer69_outs_ready
    );

  cond_br85 : entity work.cond_br_dataless(arch)
    port map(
      condition => buffer70_outs,
      condition_valid => buffer70_outs_valid,
      condition_ready => buffer70_outs_ready,
      data_valid => cond_br84_falseOut_valid,
      data_ready => cond_br84_falseOut_ready,
      clk => clk,
      rst => rst,
      trueOut_valid => cond_br85_trueOut_valid,
      trueOut_ready => cond_br85_trueOut_ready,
      falseOut_valid => cond_br85_falseOut_valid,
      falseOut_ready => cond_br85_falseOut_ready
    );

  buffer70 : entity work.tfifo(arch) generic map(1, 1)
    port map(
      ins => fork27_outs_3,
      ins_valid => fork27_outs_3_valid,
      ins_ready => fork27_outs_3_ready,
      clk => clk,
      rst => rst,
      outs => buffer70_outs,
      outs_valid => buffer70_outs_valid,
      outs_ready => buffer70_outs_ready
    );

  cond_br86 : entity work.cond_br_dataless(arch)
    port map(
      condition => buffer71_outs,
      condition_valid => buffer71_outs_valid,
      condition_ready => buffer71_outs_ready,
      data_valid => fork9_outs_0_valid,
      data_ready => fork9_outs_0_ready,
      clk => clk,
      rst => rst,
      trueOut_valid => cond_br86_trueOut_valid,
      trueOut_ready => cond_br86_trueOut_ready,
      falseOut_valid => cond_br86_falseOut_valid,
      falseOut_ready => cond_br86_falseOut_ready
    );

  buffer71 : entity work.tfifo(arch) generic map(1, 1)
    port map(
      ins => fork27_outs_2,
      ins_valid => fork27_outs_2_valid,
      ins_ready => fork27_outs_2_ready,
      clk => clk,
      rst => rst,
      outs => buffer71_outs,
      outs_valid => buffer71_outs_valid,
      outs_ready => buffer71_outs_ready
    );

  sink2 : entity work.sink_dataless(arch)
    port map(
      ins_valid => cond_br86_trueOut_valid,
      ins_ready => cond_br86_trueOut_ready,
      clk => clk,
      rst => rst
    );

  extsi45 : entity work.extsi(arch) generic map(5, 6)
    port map(
      ins => cond_br10_falseOut,
      ins_valid => cond_br10_falseOut_valid,
      ins_ready => cond_br10_falseOut_ready,
      clk => clk,
      rst => rst,
      outs => extsi45_outs,
      outs_valid => extsi45_outs_valid,
      outs_ready => extsi45_outs_ready
    );

  source5 : entity work.source(arch)
    port map(
      clk => clk,
      rst => rst,
      outs_valid => source5_outs_valid,
      outs_ready => source5_outs_ready
    );

  constant39 : entity work.handshake_constant_3(arch) generic map(5)
    port map(
      ctrl_valid => source5_outs_valid,
      ctrl_ready => source5_outs_ready,
      clk => clk,
      rst => rst,
      outs => constant39_outs,
      outs_valid => constant39_outs_valid,
      outs_ready => constant39_outs_ready
    );

  extsi46 : entity work.extsi(arch) generic map(5, 6)
    port map(
      ins => constant39_outs,
      ins_valid => constant39_outs_valid,
      ins_ready => constant39_outs_ready,
      clk => clk,
      rst => rst,
      outs => extsi46_outs,
      outs_valid => extsi46_outs_valid,
      outs_ready => extsi46_outs_ready
    );

  source6 : entity work.source(arch)
    port map(
      clk => clk,
      rst => rst,
      outs_valid => source6_outs_valid,
      outs_ready => source6_outs_ready
    );

  constant40 : entity work.handshake_constant_1(arch) generic map(2)
    port map(
      ctrl_valid => source6_outs_valid,
      ctrl_ready => source6_outs_ready,
      clk => clk,
      rst => rst,
      outs => constant40_outs,
      outs_valid => constant40_outs_valid,
      outs_ready => constant40_outs_ready
    );

  extsi47 : entity work.extsi(arch) generic map(2, 6)
    port map(
      ins => constant40_outs,
      ins_valid => constant40_outs_valid,
      ins_ready => constant40_outs_ready,
      clk => clk,
      rst => rst,
      outs => extsi47_outs,
      outs_valid => extsi47_outs_valid,
      outs_ready => extsi47_outs_ready
    );

  addi14 : entity work.addi(arch) generic map(6)
    port map(
      lhs => extsi45_outs,
      lhs_valid => extsi45_outs_valid,
      lhs_ready => extsi45_outs_ready,
      rhs => extsi47_outs,
      rhs_valid => extsi47_outs_valid,
      rhs_ready => extsi47_outs_ready,
      clk => clk,
      rst => rst,
      result => addi14_result,
      result_valid => addi14_result_valid,
      result_ready => addi14_result_ready
    );

  buffer106 : entity work.oehb(arch) generic map(6)
    port map(
      ins => addi14_result,
      ins_valid => addi14_result_valid,
      ins_ready => addi14_result_ready,
      clk => clk,
      rst => rst,
      outs => buffer106_outs,
      outs_valid => buffer106_outs_valid,
      outs_ready => buffer106_outs_ready
    );

  fork26 : entity work.handshake_fork(arch) generic map(2, 6)
    port map(
      ins => buffer106_outs,
      ins_valid => buffer106_outs_valid,
      ins_ready => buffer106_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork26_outs_0,
      outs(1) => fork26_outs_1,
      outs_valid(0) => fork26_outs_0_valid,
      outs_valid(1) => fork26_outs_1_valid,
      outs_ready(0) => fork26_outs_0_ready,
      outs_ready(1) => fork26_outs_1_ready
    );

  trunci9 : entity work.trunci(arch) generic map(6, 5)
    port map(
      ins => fork26_outs_0,
      ins_valid => fork26_outs_0_valid,
      ins_ready => fork26_outs_0_ready,
      clk => clk,
      rst => rst,
      outs => trunci9_outs,
      outs_valid => trunci9_outs_valid,
      outs_ready => trunci9_outs_ready
    );

  cmpi1 : entity work.handshake_cmpi_0(arch) generic map(6)
    port map(
      lhs => fork26_outs_1,
      lhs_valid => fork26_outs_1_valid,
      lhs_ready => fork26_outs_1_ready,
      rhs => extsi46_outs,
      rhs_valid => extsi46_outs_valid,
      rhs_ready => extsi46_outs_ready,
      clk => clk,
      rst => rst,
      result => cmpi1_result,
      result_valid => cmpi1_result_valid,
      result_ready => cmpi1_result_ready
    );

  buffer107 : entity work.oehb(arch) generic map(1)
    port map(
      ins => cmpi1_result,
      ins_valid => cmpi1_result_valid,
      ins_ready => cmpi1_result_ready,
      clk => clk,
      rst => rst,
      outs => buffer107_outs,
      outs_valid => buffer107_outs_valid,
      outs_ready => buffer107_outs_ready
    );

  fork27 : entity work.handshake_fork(arch) generic map(8, 1)
    port map(
      ins => buffer107_outs,
      ins_valid => buffer107_outs_valid,
      ins_ready => buffer107_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork27_outs_0,
      outs(1) => fork27_outs_1,
      outs(2) => fork27_outs_2,
      outs(3) => fork27_outs_3,
      outs(4) => fork27_outs_4,
      outs(5) => fork27_outs_5,
      outs(6) => fork27_outs_6,
      outs(7) => fork27_outs_7,
      outs_valid(0) => fork27_outs_0_valid,
      outs_valid(1) => fork27_outs_1_valid,
      outs_valid(2) => fork27_outs_2_valid,
      outs_valid(3) => fork27_outs_3_valid,
      outs_valid(4) => fork27_outs_4_valid,
      outs_valid(5) => fork27_outs_5_valid,
      outs_valid(6) => fork27_outs_6_valid,
      outs_valid(7) => fork27_outs_7_valid,
      outs_ready(0) => fork27_outs_0_ready,
      outs_ready(1) => fork27_outs_1_ready,
      outs_ready(2) => fork27_outs_2_ready,
      outs_ready(3) => fork27_outs_3_ready,
      outs_ready(4) => fork27_outs_4_ready,
      outs_ready(5) => fork27_outs_5_ready,
      outs_ready(6) => fork27_outs_6_ready,
      outs_ready(7) => fork27_outs_7_ready
    );

  cond_br12 : entity work.cond_br(arch) generic map(5)
    port map(
      condition => fork27_outs_0,
      condition_valid => fork27_outs_0_valid,
      condition_ready => fork27_outs_0_ready,
      data => trunci9_outs,
      data_valid => trunci9_outs_valid,
      data_ready => trunci9_outs_ready,
      clk => clk,
      rst => rst,
      trueOut => cond_br12_trueOut,
      trueOut_valid => cond_br12_trueOut_valid,
      trueOut_ready => cond_br12_trueOut_ready,
      falseOut => cond_br12_falseOut,
      falseOut_valid => cond_br12_falseOut_valid,
      falseOut_ready => cond_br12_falseOut_ready
    );

  sink4 : entity work.sink(arch) generic map(5)
    port map(
      ins => cond_br12_falseOut,
      ins_valid => cond_br12_falseOut_valid,
      ins_ready => cond_br12_falseOut_ready,
      clk => clk,
      rst => rst
    );

  buffer104 : entity work.oehb(arch) generic map(32)
    port map(
      ins => cond_br7_falseOut,
      ins_valid => cond_br7_falseOut_valid,
      ins_ready => cond_br7_falseOut_ready,
      clk => clk,
      rst => rst,
      outs => buffer104_outs,
      outs_valid => buffer104_outs_valid,
      outs_ready => buffer104_outs_ready
    );

  cond_br13 : entity work.cond_br(arch) generic map(32)
    port map(
      condition => buffer75_outs,
      condition_valid => buffer75_outs_valid,
      condition_ready => buffer75_outs_ready,
      data => buffer104_outs,
      data_valid => buffer104_outs_valid,
      data_ready => buffer104_outs_ready,
      clk => clk,
      rst => rst,
      trueOut => cond_br13_trueOut,
      trueOut_valid => cond_br13_trueOut_valid,
      trueOut_ready => cond_br13_trueOut_ready,
      falseOut => cond_br13_falseOut,
      falseOut_valid => cond_br13_falseOut_valid,
      falseOut_ready => cond_br13_falseOut_ready
    );

  buffer75 : entity work.tfifo(arch) generic map(1, 1)
    port map(
      ins => fork27_outs_5,
      ins_valid => fork27_outs_5_valid,
      ins_ready => fork27_outs_5_ready,
      clk => clk,
      rst => rst,
      outs => buffer75_outs,
      outs_valid => buffer75_outs_valid,
      outs_ready => buffer75_outs_ready
    );

  buffer105 : entity work.oehb(arch) generic map(32)
    port map(
      ins => cond_br8_falseOut,
      ins_valid => cond_br8_falseOut_valid,
      ins_ready => cond_br8_falseOut_ready,
      clk => clk,
      rst => rst,
      outs => buffer105_outs,
      outs_valid => buffer105_outs_valid,
      outs_ready => buffer105_outs_ready
    );

  cond_br14 : entity work.cond_br(arch) generic map(32)
    port map(
      condition => buffer76_outs,
      condition_valid => buffer76_outs_valid,
      condition_ready => buffer76_outs_ready,
      data => buffer105_outs,
      data_valid => buffer105_outs_valid,
      data_ready => buffer105_outs_ready,
      clk => clk,
      rst => rst,
      trueOut => cond_br14_trueOut,
      trueOut_valid => cond_br14_trueOut_valid,
      trueOut_ready => cond_br14_trueOut_ready,
      falseOut => cond_br14_falseOut,
      falseOut_valid => cond_br14_falseOut_valid,
      falseOut_ready => cond_br14_falseOut_ready
    );

  buffer76 : entity work.tfifo(arch) generic map(1, 1)
    port map(
      ins => fork27_outs_6,
      ins_valid => fork27_outs_6_valid,
      ins_ready => fork27_outs_6_ready,
      clk => clk,
      rst => rst,
      outs => buffer76_outs,
      outs_valid => buffer76_outs_valid,
      outs_ready => buffer76_outs_ready
    );

  cond_br15 : entity work.cond_br(arch) generic map(5)
    port map(
      condition => fork27_outs_1,
      condition_valid => fork27_outs_1_valid,
      condition_ready => fork27_outs_1_ready,
      data => cond_br9_falseOut,
      data_valid => cond_br9_falseOut_valid,
      data_ready => cond_br9_falseOut_ready,
      clk => clk,
      rst => rst,
      trueOut => cond_br15_trueOut,
      trueOut_valid => cond_br15_trueOut_valid,
      trueOut_ready => cond_br15_trueOut_ready,
      falseOut => cond_br15_falseOut,
      falseOut_valid => cond_br15_falseOut_valid,
      falseOut_ready => cond_br15_falseOut_ready
    );

  cond_br16 : entity work.cond_br_dataless(arch)
    port map(
      condition => buffer78_outs,
      condition_valid => buffer78_outs_valid,
      condition_ready => buffer78_outs_ready,
      data_valid => cond_br11_falseOut_valid,
      data_ready => cond_br11_falseOut_ready,
      clk => clk,
      rst => rst,
      trueOut_valid => cond_br16_trueOut_valid,
      trueOut_ready => cond_br16_trueOut_ready,
      falseOut_valid => cond_br16_falseOut_valid,
      falseOut_ready => cond_br16_falseOut_ready
    );

  buffer78 : entity work.tfifo(arch) generic map(1, 1)
    port map(
      ins => fork27_outs_7,
      ins_valid => fork27_outs_7_valid,
      ins_ready => fork27_outs_7_ready,
      clk => clk,
      rst => rst,
      outs => buffer78_outs,
      outs_valid => buffer78_outs_valid,
      outs_ready => buffer78_outs_ready
    );

  cond_br87 : entity work.cond_br_dataless(arch)
    port map(
      condition => fork30_outs_2,
      condition_valid => fork30_outs_2_valid,
      condition_ready => fork30_outs_2_ready,
      data_valid => cond_br86_falseOut_valid,
      data_ready => cond_br86_falseOut_ready,
      clk => clk,
      rst => rst,
      trueOut_valid => cond_br87_trueOut_valid,
      trueOut_ready => cond_br87_trueOut_ready,
      falseOut_valid => cond_br87_falseOut_valid,
      falseOut_ready => cond_br87_falseOut_ready
    );

  sink5 : entity work.sink_dataless(arch)
    port map(
      ins_valid => cond_br87_trueOut_valid,
      ins_ready => cond_br87_trueOut_ready,
      clk => clk,
      rst => rst
    );

  cond_br88 : entity work.cond_br_dataless(arch)
    port map(
      condition => buffer80_outs,
      condition_valid => buffer80_outs_valid,
      condition_ready => buffer80_outs_ready,
      data_valid => cond_br85_falseOut_valid,
      data_ready => cond_br85_falseOut_ready,
      clk => clk,
      rst => rst,
      trueOut_valid => cond_br88_trueOut_valid,
      trueOut_ready => cond_br88_trueOut_ready,
      falseOut_valid => cond_br88_falseOut_valid,
      falseOut_ready => cond_br88_falseOut_ready
    );

  buffer80 : entity work.tfifo(arch) generic map(1, 1)
    port map(
      ins => fork30_outs_1,
      ins_valid => fork30_outs_1_valid,
      ins_ready => fork30_outs_1_ready,
      clk => clk,
      rst => rst,
      outs => buffer80_outs,
      outs_valid => buffer80_outs_valid,
      outs_ready => buffer80_outs_ready
    );

  buffer108 : entity work.oehb(arch) generic map(5)
    port map(
      ins => cond_br15_falseOut,
      ins_valid => cond_br15_falseOut_valid,
      ins_ready => cond_br15_falseOut_ready,
      clk => clk,
      rst => rst,
      outs => buffer108_outs,
      outs_valid => buffer108_outs_valid,
      outs_ready => buffer108_outs_ready
    );

  extsi48 : entity work.extsi(arch) generic map(5, 6)
    port map(
      ins => buffer108_outs,
      ins_valid => buffer108_outs_valid,
      ins_ready => buffer108_outs_ready,
      clk => clk,
      rst => rst,
      outs => extsi48_outs,
      outs_valid => extsi48_outs_valid,
      outs_ready => extsi48_outs_ready
    );

  fork28 : entity work.fork_dataless(arch) generic map(2)
    port map(
      ins_valid => cond_br16_falseOut_valid,
      ins_ready => cond_br16_falseOut_ready,
      clk => clk,
      rst => rst,
      outs_valid(0) => fork28_outs_0_valid,
      outs_valid(1) => fork28_outs_1_valid,
      outs_ready(0) => fork28_outs_0_ready,
      outs_ready(1) => fork28_outs_1_ready
    );

  constant41 : entity work.handshake_constant_0(arch) generic map(1)
    port map(
      ctrl_valid => fork28_outs_0_valid,
      ctrl_ready => fork28_outs_0_ready,
      clk => clk,
      rst => rst,
      outs => constant41_outs,
      outs_valid => constant41_outs_valid,
      outs_ready => constant41_outs_ready
    );

  source7 : entity work.source(arch)
    port map(
      clk => clk,
      rst => rst,
      outs_valid => source7_outs_valid,
      outs_ready => source7_outs_ready
    );

  constant42 : entity work.handshake_constant_3(arch) generic map(5)
    port map(
      ctrl_valid => source7_outs_valid,
      ctrl_ready => source7_outs_ready,
      clk => clk,
      rst => rst,
      outs => constant42_outs,
      outs_valid => constant42_outs_valid,
      outs_ready => constant42_outs_ready
    );

  extsi49 : entity work.extsi(arch) generic map(5, 6)
    port map(
      ins => constant42_outs,
      ins_valid => constant42_outs_valid,
      ins_ready => constant42_outs_ready,
      clk => clk,
      rst => rst,
      outs => extsi49_outs,
      outs_valid => extsi49_outs_valid,
      outs_ready => extsi49_outs_ready
    );

  source8 : entity work.source(arch)
    port map(
      clk => clk,
      rst => rst,
      outs_valid => source8_outs_valid,
      outs_ready => source8_outs_ready
    );

  constant43 : entity work.handshake_constant_1(arch) generic map(2)
    port map(
      ctrl_valid => source8_outs_valid,
      ctrl_ready => source8_outs_ready,
      clk => clk,
      rst => rst,
      outs => constant43_outs,
      outs_valid => constant43_outs_valid,
      outs_ready => constant43_outs_ready
    );

  extsi50 : entity work.extsi(arch) generic map(2, 6)
    port map(
      ins => constant43_outs,
      ins_valid => constant43_outs_valid,
      ins_ready => constant43_outs_ready,
      clk => clk,
      rst => rst,
      outs => extsi50_outs,
      outs_valid => extsi50_outs_valid,
      outs_ready => extsi50_outs_ready
    );

  addi15 : entity work.addi(arch) generic map(6)
    port map(
      lhs => extsi48_outs,
      lhs_valid => extsi48_outs_valid,
      lhs_ready => extsi48_outs_ready,
      rhs => extsi50_outs,
      rhs_valid => extsi50_outs_valid,
      rhs_ready => extsi50_outs_ready,
      clk => clk,
      rst => rst,
      result => addi15_result,
      result_valid => addi15_result_valid,
      result_ready => addi15_result_ready
    );

  buffer109 : entity work.oehb(arch) generic map(6)
    port map(
      ins => addi15_result,
      ins_valid => addi15_result_valid,
      ins_ready => addi15_result_ready,
      clk => clk,
      rst => rst,
      outs => buffer109_outs,
      outs_valid => buffer109_outs_valid,
      outs_ready => buffer109_outs_ready
    );

  fork29 : entity work.handshake_fork(arch) generic map(2, 6)
    port map(
      ins => buffer109_outs,
      ins_valid => buffer109_outs_valid,
      ins_ready => buffer109_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork29_outs_0,
      outs(1) => fork29_outs_1,
      outs_valid(0) => fork29_outs_0_valid,
      outs_valid(1) => fork29_outs_1_valid,
      outs_ready(0) => fork29_outs_0_ready,
      outs_ready(1) => fork29_outs_1_ready
    );

  trunci10 : entity work.trunci(arch) generic map(6, 5)
    port map(
      ins => fork29_outs_0,
      ins_valid => fork29_outs_0_valid,
      ins_ready => fork29_outs_0_ready,
      clk => clk,
      rst => rst,
      outs => trunci10_outs,
      outs_valid => trunci10_outs_valid,
      outs_ready => trunci10_outs_ready
    );

  cmpi2 : entity work.handshake_cmpi_0(arch) generic map(6)
    port map(
      lhs => fork29_outs_1,
      lhs_valid => fork29_outs_1_valid,
      lhs_ready => fork29_outs_1_ready,
      rhs => extsi49_outs,
      rhs_valid => extsi49_outs_valid,
      rhs_ready => extsi49_outs_ready,
      clk => clk,
      rst => rst,
      result => cmpi2_result,
      result_valid => cmpi2_result_valid,
      result_ready => cmpi2_result_ready
    );

  buffer114 : entity work.oehb(arch) generic map(1)
    port map(
      ins => cmpi2_result,
      ins_valid => cmpi2_result_valid,
      ins_ready => cmpi2_result_ready,
      clk => clk,
      rst => rst,
      outs => buffer114_outs,
      outs_valid => buffer114_outs_valid,
      outs_ready => buffer114_outs_ready
    );

  fork30 : entity work.handshake_fork(arch) generic map(8, 1)
    port map(
      ins => buffer114_outs,
      ins_valid => buffer114_outs_valid,
      ins_ready => buffer114_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork30_outs_0,
      outs(1) => fork30_outs_1,
      outs(2) => fork30_outs_2,
      outs(3) => fork30_outs_3,
      outs(4) => fork30_outs_4,
      outs(5) => fork30_outs_5,
      outs(6) => fork30_outs_6,
      outs(7) => fork30_outs_7,
      outs_valid(0) => fork30_outs_0_valid,
      outs_valid(1) => fork30_outs_1_valid,
      outs_valid(2) => fork30_outs_2_valid,
      outs_valid(3) => fork30_outs_3_valid,
      outs_valid(4) => fork30_outs_4_valid,
      outs_valid(5) => fork30_outs_5_valid,
      outs_valid(6) => fork30_outs_6_valid,
      outs_valid(7) => fork30_outs_7_valid,
      outs_ready(0) => fork30_outs_0_ready,
      outs_ready(1) => fork30_outs_1_ready,
      outs_ready(2) => fork30_outs_2_ready,
      outs_ready(3) => fork30_outs_3_ready,
      outs_ready(4) => fork30_outs_4_ready,
      outs_ready(5) => fork30_outs_5_ready,
      outs_ready(6) => fork30_outs_6_ready,
      outs_ready(7) => fork30_outs_7_ready
    );

  cond_br17 : entity work.cond_br(arch) generic map(5)
    port map(
      condition => fork30_outs_0,
      condition_valid => fork30_outs_0_valid,
      condition_ready => fork30_outs_0_ready,
      data => trunci10_outs,
      data_valid => trunci10_outs_valid,
      data_ready => trunci10_outs_ready,
      clk => clk,
      rst => rst,
      trueOut => cond_br17_trueOut,
      trueOut_valid => cond_br17_trueOut_valid,
      trueOut_ready => cond_br17_trueOut_ready,
      falseOut => cond_br17_falseOut,
      falseOut_valid => cond_br17_falseOut_valid,
      falseOut_ready => cond_br17_falseOut_ready
    );

  sink7 : entity work.sink(arch) generic map(5)
    port map(
      ins => cond_br17_falseOut,
      ins_valid => cond_br17_falseOut_valid,
      ins_ready => cond_br17_falseOut_ready,
      clk => clk,
      rst => rst
    );

  cond_br18 : entity work.cond_br(arch) generic map(32)
    port map(
      condition => fork30_outs_4,
      condition_valid => fork30_outs_4_valid,
      condition_ready => fork30_outs_4_ready,
      data => cond_br13_falseOut,
      data_valid => cond_br13_falseOut_valid,
      data_ready => cond_br13_falseOut_ready,
      clk => clk,
      rst => rst,
      trueOut => cond_br18_trueOut,
      trueOut_valid => cond_br18_trueOut_valid,
      trueOut_ready => cond_br18_trueOut_ready,
      falseOut => cond_br18_falseOut,
      falseOut_valid => cond_br18_falseOut_valid,
      falseOut_ready => cond_br18_falseOut_ready
    );

  sink8 : entity work.sink(arch) generic map(32)
    port map(
      ins => cond_br18_falseOut,
      ins_valid => cond_br18_falseOut_valid,
      ins_ready => cond_br18_falseOut_ready,
      clk => clk,
      rst => rst
    );

  cond_br19 : entity work.cond_br(arch) generic map(32)
    port map(
      condition => fork30_outs_5,
      condition_valid => fork30_outs_5_valid,
      condition_ready => fork30_outs_5_ready,
      data => cond_br14_falseOut,
      data_valid => cond_br14_falseOut_valid,
      data_ready => cond_br14_falseOut_ready,
      clk => clk,
      rst => rst,
      trueOut => cond_br19_trueOut,
      trueOut_valid => cond_br19_trueOut_valid,
      trueOut_ready => cond_br19_trueOut_ready,
      falseOut => cond_br19_falseOut,
      falseOut_valid => cond_br19_falseOut_valid,
      falseOut_ready => cond_br19_falseOut_ready
    );

  cond_br20 : entity work.cond_br_dataless(arch)
    port map(
      condition => fork30_outs_6,
      condition_valid => fork30_outs_6_valid,
      condition_ready => fork30_outs_6_ready,
      data_valid => fork28_outs_1_valid,
      data_ready => fork28_outs_1_ready,
      clk => clk,
      rst => rst,
      trueOut_valid => cond_br20_trueOut_valid,
      trueOut_ready => cond_br20_trueOut_ready,
      falseOut_valid => cond_br20_falseOut_valid,
      falseOut_ready => cond_br20_falseOut_ready
    );

  cond_br21 : entity work.cond_br(arch) generic map(1)
    port map(
      condition => fork30_outs_7,
      condition_valid => fork30_outs_7_valid,
      condition_ready => fork30_outs_7_ready,
      data => constant41_outs,
      data_valid => constant41_outs_valid,
      data_ready => constant41_outs_ready,
      clk => clk,
      rst => rst,
      trueOut => cond_br21_trueOut,
      trueOut_valid => cond_br21_trueOut_valid,
      trueOut_ready => cond_br21_trueOut_ready,
      falseOut => cond_br21_falseOut,
      falseOut_valid => cond_br21_falseOut_valid,
      falseOut_ready => cond_br21_falseOut_ready
    );

  sink9 : entity work.sink(arch) generic map(1)
    port map(
      ins => cond_br21_trueOut,
      ins_valid => cond_br21_trueOut_valid,
      ins_ready => cond_br21_trueOut_ready,
      clk => clk,
      rst => rst
    );

  extsi31 : entity work.extsi(arch) generic map(1, 5)
    port map(
      ins => cond_br21_falseOut,
      ins_valid => cond_br21_falseOut_valid,
      ins_ready => cond_br21_falseOut_ready,
      clk => clk,
      rst => rst,
      outs => extsi31_outs,
      outs_valid => extsi31_outs_valid,
      outs_ready => extsi31_outs_ready
    );

  init14 : entity work.tehb_init(arch) generic map(1, 0)
    port map(
      ins => fork69_outs_4,
      ins_valid => fork69_outs_4_valid,
      ins_ready => fork69_outs_4_ready,
      clk => clk,
      rst => rst,
      outs => init14_outs,
      outs_valid => init14_outs_valid,
      outs_ready => init14_outs_ready
    );

  fork31 : entity work.handshake_fork(arch) generic map(3, 1)
    port map(
      ins => init14_outs,
      ins_valid => init14_outs_valid,
      ins_ready => init14_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork31_outs_0,
      outs(1) => fork31_outs_1,
      outs(2) => fork31_outs_2,
      outs_valid(0) => fork31_outs_0_valid,
      outs_valid(1) => fork31_outs_1_valid,
      outs_valid(2) => fork31_outs_2_valid,
      outs_ready(0) => fork31_outs_0_ready,
      outs_ready(1) => fork31_outs_1_ready,
      outs_ready(2) => fork31_outs_2_ready
    );

  buffer215 : entity work.oehb_dataless(arch)
    port map(
      ins_valid => cond_br99_trueOut_valid,
      ins_ready => cond_br99_trueOut_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer215_outs_valid,
      outs_ready => buffer215_outs_ready
    );

  mux35 : entity work.mux_dataless(arch) generic map(2, 1)
    port map(
      index => buffer89_outs,
      index_valid => buffer89_outs_valid,
      index_ready => buffer89_outs_ready,
      ins_valid(0) => cond_br88_falseOut_valid,
      ins_valid(1) => buffer215_outs_valid,
      ins_ready(0) => cond_br88_falseOut_ready,
      ins_ready(1) => buffer215_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => mux35_outs_valid,
      outs_ready => mux35_outs_ready
    );

  buffer89 : entity work.tfifo(arch) generic map(1, 1)
    port map(
      ins => fork31_outs_2,
      ins_valid => fork31_outs_2_valid,
      ins_ready => fork31_outs_2_ready,
      clk => clk,
      rst => rst,
      outs => buffer89_outs,
      outs_valid => buffer89_outs_valid,
      outs_ready => buffer89_outs_ready
    );

  buffer115 : entity work.tehb_dataless(arch)
    port map(
      ins_valid => mux35_outs_valid,
      ins_ready => mux35_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer115_outs_valid,
      outs_ready => buffer115_outs_ready
    );

  fork32 : entity work.fork_dataless(arch) generic map(2)
    port map(
      ins_valid => buffer115_outs_valid,
      ins_ready => buffer115_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid(0) => fork32_outs_0_valid,
      outs_valid(1) => fork32_outs_1_valid,
      outs_ready(0) => fork32_outs_0_ready,
      outs_ready(1) => fork32_outs_1_ready
    );

  mux36 : entity work.mux_dataless(arch) generic map(2, 1)
    port map(
      index => buffer90_outs,
      index_valid => buffer90_outs_valid,
      index_ready => buffer90_outs_ready,
      ins_valid(0) => cond_br87_falseOut_valid,
      ins_valid(1) => cond_br98_trueOut_valid,
      ins_ready(0) => cond_br87_falseOut_ready,
      ins_ready(1) => cond_br98_trueOut_ready,
      clk => clk,
      rst => rst,
      outs_valid => mux36_outs_valid,
      outs_ready => mux36_outs_ready
    );

  buffer90 : entity work.tfifo(arch) generic map(1, 1)
    port map(
      ins => fork31_outs_1,
      ins_valid => fork31_outs_1_valid,
      ins_ready => fork31_outs_1_ready,
      clk => clk,
      rst => rst,
      outs => buffer90_outs,
      outs_valid => buffer90_outs_valid,
      outs_ready => buffer90_outs_ready
    );

  buffer116 : entity work.oehb_dataless(arch)
    port map(
      ins_valid => mux36_outs_valid,
      ins_ready => mux36_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer116_outs_valid,
      outs_ready => buffer116_outs_ready
    );

  buffer117 : entity work.tehb_dataless(arch)
    port map(
      ins_valid => buffer116_outs_valid,
      ins_ready => buffer116_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer117_outs_valid,
      outs_ready => buffer117_outs_ready
    );

  fork33 : entity work.fork_dataless(arch) generic map(2)
    port map(
      ins_valid => buffer117_outs_valid,
      ins_ready => buffer117_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid(0) => fork33_outs_0_valid,
      outs_valid(1) => fork33_outs_1_valid,
      outs_ready(0) => fork33_outs_0_ready,
      outs_ready(1) => fork33_outs_1_ready
    );

  mux40 : entity work.mux_dataless(arch) generic map(2, 1)
    port map(
      index => buffer91_outs,
      index_valid => buffer91_outs_valid,
      index_ready => buffer91_outs_ready,
      ins_valid(0) => fork0_outs_2_valid,
      ins_valid(1) => cond_br97_trueOut_valid,
      ins_ready(0) => fork0_outs_2_ready,
      ins_ready(1) => cond_br97_trueOut_ready,
      clk => clk,
      rst => rst,
      outs_valid => mux40_outs_valid,
      outs_ready => mux40_outs_ready
    );

  buffer91 : entity work.tfifo(arch) generic map(1, 1)
    port map(
      ins => fork31_outs_0,
      ins_valid => fork31_outs_0_valid,
      ins_ready => fork31_outs_0_ready,
      clk => clk,
      rst => rst,
      outs => buffer91_outs,
      outs_valid => buffer91_outs_valid,
      outs_ready => buffer91_outs_ready
    );

  mux12 : entity work.mux(arch) generic map(2, 5, 1)
    port map(
      index => fork34_outs_0,
      index_valid => fork34_outs_0_valid,
      index_ready => fork34_outs_0_ready,
      ins(0) => extsi31_outs,
      ins(1) => cond_br31_trueOut,
      ins_valid(0) => extsi31_outs_valid,
      ins_valid(1) => cond_br31_trueOut_valid,
      ins_ready(0) => extsi31_outs_ready,
      ins_ready(1) => cond_br31_trueOut_ready,
      clk => clk,
      rst => rst,
      outs => mux12_outs,
      outs_valid => mux12_outs_valid,
      outs_ready => mux12_outs_ready
    );

  mux13 : entity work.mux(arch) generic map(2, 32, 1)
    port map(
      index => fork34_outs_1,
      index_valid => fork34_outs_1_valid,
      index_ready => fork34_outs_1_ready,
      ins(0) => cond_br19_falseOut,
      ins(1) => cond_br32_trueOut,
      ins_valid(0) => cond_br19_falseOut_valid,
      ins_valid(1) => cond_br32_trueOut_valid,
      ins_ready(0) => cond_br19_falseOut_ready,
      ins_ready(1) => cond_br32_trueOut_ready,
      clk => clk,
      rst => rst,
      outs => mux13_outs,
      outs_valid => mux13_outs_valid,
      outs_ready => mux13_outs_ready
    );

  control_merge5 : entity work.control_merge_dataless(arch) generic map(2, 1)
    port map(
      ins_valid(0) => cond_br20_falseOut_valid,
      ins_valid(1) => cond_br33_trueOut_valid,
      ins_ready(0) => cond_br20_falseOut_ready,
      ins_ready(1) => cond_br33_trueOut_ready,
      clk => clk,
      rst => rst,
      outs_valid => control_merge5_outs_valid,
      outs_ready => control_merge5_outs_ready,
      index => control_merge5_index,
      index_valid => control_merge5_index_valid,
      index_ready => control_merge5_index_ready
    );

  fork34 : entity work.handshake_fork(arch) generic map(2, 1)
    port map(
      ins => control_merge5_index,
      ins_valid => control_merge5_index_valid,
      ins_ready => control_merge5_index_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork34_outs_0,
      outs(1) => fork34_outs_1,
      outs_valid(0) => fork34_outs_0_valid,
      outs_valid(1) => fork34_outs_1_valid,
      outs_ready(0) => fork34_outs_0_ready,
      outs_ready(1) => fork34_outs_1_ready
    );

  fork35 : entity work.fork_dataless(arch) generic map(2)
    port map(
      ins_valid => control_merge5_outs_valid,
      ins_ready => control_merge5_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid(0) => fork35_outs_0_valid,
      outs_valid(1) => fork35_outs_1_valid,
      outs_ready(0) => fork35_outs_0_ready,
      outs_ready(1) => fork35_outs_1_ready
    );

  constant44 : entity work.handshake_constant_0(arch) generic map(1)
    port map(
      ctrl_valid => fork35_outs_0_valid,
      ctrl_ready => fork35_outs_0_ready,
      clk => clk,
      rst => rst,
      outs => constant44_outs,
      outs_valid => constant44_outs_valid,
      outs_ready => constant44_outs_ready
    );

  extsi30 : entity work.extsi(arch) generic map(1, 5)
    port map(
      ins => constant44_outs,
      ins_valid => constant44_outs_valid,
      ins_ready => constant44_outs_ready,
      clk => clk,
      rst => rst,
      outs => extsi30_outs,
      outs_valid => extsi30_outs_valid,
      outs_ready => extsi30_outs_ready
    );

  buffer129 : entity work.oehb(arch) generic map(32)
    port map(
      ins => mux13_outs,
      ins_valid => mux13_outs_valid,
      ins_ready => mux13_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer129_outs,
      outs_valid => buffer129_outs_valid,
      outs_ready => buffer129_outs_ready
    );

  buffer130 : entity work.tehb(arch) generic map(32)
    port map(
      ins => buffer129_outs,
      ins_valid => buffer129_outs_valid,
      ins_ready => buffer129_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer130_outs,
      outs_valid => buffer130_outs_valid,
      outs_ready => buffer130_outs_ready
    );

  buffer123 : entity work.tehb(arch) generic map(5)
    port map(
      ins => mux12_outs,
      ins_valid => mux12_outs_valid,
      ins_ready => mux12_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer123_outs,
      outs_valid => buffer123_outs_valid,
      outs_ready => buffer123_outs_ready
    );

  init20 : entity work.tehb_init(arch) generic map(1, 0)
    port map(
      ins => fork67_outs_5,
      ins_valid => fork67_outs_5_valid,
      ins_ready => fork67_outs_5_ready,
      clk => clk,
      rst => rst,
      outs => init20_outs,
      outs_valid => init20_outs_valid,
      outs_ready => init20_outs_ready
    );

  fork36 : entity work.handshake_fork(arch) generic map(3, 1)
    port map(
      ins => init20_outs,
      ins_valid => init20_outs_valid,
      ins_ready => init20_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork36_outs_0,
      outs(1) => fork36_outs_1,
      outs(2) => fork36_outs_2,
      outs_valid(0) => fork36_outs_0_valid,
      outs_valid(1) => fork36_outs_1_valid,
      outs_valid(2) => fork36_outs_2_valid,
      outs_ready(0) => fork36_outs_0_ready,
      outs_ready(1) => fork36_outs_1_ready,
      outs_ready(2) => fork36_outs_2_ready
    );

  mux41 : entity work.mux_dataless(arch) generic map(2, 1)
    port map(
      index => buffer95_outs,
      index_valid => buffer95_outs_valid,
      index_ready => buffer95_outs_ready,
      ins_valid(0) => fork32_outs_1_valid,
      ins_valid(1) => cond_br95_trueOut_valid,
      ins_ready(0) => fork32_outs_1_ready,
      ins_ready(1) => cond_br95_trueOut_ready,
      clk => clk,
      rst => rst,
      outs_valid => mux41_outs_valid,
      outs_ready => mux41_outs_ready
    );

  buffer95 : entity work.tfifo(arch) generic map(1, 1)
    port map(
      ins => fork36_outs_2,
      ins_valid => fork36_outs_2_valid,
      ins_ready => fork36_outs_2_ready,
      clk => clk,
      rst => rst,
      outs => buffer95_outs,
      outs_valid => buffer95_outs_valid,
      outs_ready => buffer95_outs_ready
    );

  buffer131 : entity work.oehb_dataless(arch)
    port map(
      ins_valid => mux41_outs_valid,
      ins_ready => mux41_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer131_outs_valid,
      outs_ready => buffer131_outs_ready
    );

  buffer132 : entity work.tehb_dataless(arch)
    port map(
      ins_valid => buffer131_outs_valid,
      ins_ready => buffer131_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer132_outs_valid,
      outs_ready => buffer132_outs_ready
    );

  fork37 : entity work.fork_dataless(arch) generic map(2)
    port map(
      ins_valid => buffer132_outs_valid,
      ins_ready => buffer132_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid(0) => fork37_outs_0_valid,
      outs_valid(1) => fork37_outs_1_valid,
      outs_ready(0) => fork37_outs_0_ready,
      outs_ready(1) => fork37_outs_1_ready
    );

  mux42 : entity work.mux_dataless(arch) generic map(2, 1)
    port map(
      index => buffer96_outs,
      index_valid => buffer96_outs_valid,
      index_ready => buffer96_outs_ready,
      ins_valid(0) => fork33_outs_1_valid,
      ins_valid(1) => cond_br94_trueOut_valid,
      ins_ready(0) => fork33_outs_1_ready,
      ins_ready(1) => cond_br94_trueOut_ready,
      clk => clk,
      rst => rst,
      outs_valid => mux42_outs_valid,
      outs_ready => mux42_outs_ready
    );

  buffer96 : entity work.tfifo(arch) generic map(1, 1)
    port map(
      ins => fork36_outs_1,
      ins_valid => fork36_outs_1_valid,
      ins_ready => fork36_outs_1_ready,
      clk => clk,
      rst => rst,
      outs => buffer96_outs,
      outs_valid => buffer96_outs_valid,
      outs_ready => buffer96_outs_ready
    );

  buffer133 : entity work.oehb_dataless(arch)
    port map(
      ins_valid => mux42_outs_valid,
      ins_ready => mux42_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer133_outs_valid,
      outs_ready => buffer133_outs_ready
    );

  buffer135 : entity work.tehb_dataless(arch)
    port map(
      ins_valid => buffer133_outs_valid,
      ins_ready => buffer133_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer135_outs_valid,
      outs_ready => buffer135_outs_ready
    );

  fork38 : entity work.fork_dataless(arch) generic map(2)
    port map(
      ins_valid => buffer135_outs_valid,
      ins_ready => buffer135_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid(0) => fork38_outs_0_valid,
      outs_valid(1) => fork38_outs_1_valid,
      outs_ready(0) => fork38_outs_0_ready,
      outs_ready(1) => fork38_outs_1_ready
    );

  buffer121 : entity work.tehb_dataless(arch)
    port map(
      ins_valid => mux40_outs_valid,
      ins_ready => mux40_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer121_outs_valid,
      outs_ready => buffer121_outs_ready
    );

  mux46 : entity work.mux_dataless(arch) generic map(2, 1)
    port map(
      index => buffer97_outs,
      index_valid => buffer97_outs_valid,
      index_ready => buffer97_outs_ready,
      ins_valid(0) => buffer121_outs_valid,
      ins_valid(1) => cond_br96_trueOut_valid,
      ins_ready(0) => buffer121_outs_ready,
      ins_ready(1) => cond_br96_trueOut_ready,
      clk => clk,
      rst => rst,
      outs_valid => mux46_outs_valid,
      outs_ready => mux46_outs_ready
    );

  buffer97 : entity work.tfifo(arch) generic map(1, 1)
    port map(
      ins => fork36_outs_0,
      ins_valid => fork36_outs_0_valid,
      ins_ready => fork36_outs_0_ready,
      clk => clk,
      rst => rst,
      outs => buffer97_outs,
      outs_valid => buffer97_outs_valid,
      outs_ready => buffer97_outs_ready
    );

  unbundle2 : entity work.unbundle(arch) generic map(32)
    port map(
      ins => buffer98_outs,
      ins_valid => buffer98_outs_valid,
      ins_ready => buffer98_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => unbundle2_outs_0_valid,
      outs_ready => unbundle2_outs_0_ready,
      outs => unbundle2_outs_1
    );

  buffer98 : entity work.tfifo(arch) generic map(1, 32)
    port map(
      ins => fork47_outs_0,
      ins_valid => fork47_outs_0_valid,
      ins_ready => fork47_outs_0_ready,
      clk => clk,
      rst => rst,
      outs => buffer98_outs,
      outs_valid => buffer98_outs_valid,
      outs_ready => buffer98_outs_ready
    );

  mux14 : entity work.mux(arch) generic map(2, 5, 1)
    port map(
      index => fork43_outs_1,
      index_valid => fork43_outs_1_valid,
      index_ready => fork43_outs_1_ready,
      ins(0) => extsi30_outs,
      ins(1) => cond_br27_trueOut,
      ins_valid(0) => extsi30_outs_valid,
      ins_valid(1) => cond_br27_trueOut_valid,
      ins_ready(0) => extsi30_outs_ready,
      ins_ready(1) => cond_br27_trueOut_ready,
      clk => clk,
      rst => rst,
      outs => mux14_outs,
      outs_valid => mux14_outs_valid,
      outs_ready => mux14_outs_ready
    );

  buffer142 : entity work.tehb(arch) generic map(5)
    port map(
      ins => mux14_outs,
      ins_valid => mux14_outs_valid,
      ins_ready => mux14_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer142_outs,
      outs_valid => buffer142_outs_valid,
      outs_ready => buffer142_outs_ready
    );

  fork39 : entity work.handshake_fork(arch) generic map(3, 5)
    port map(
      ins => buffer142_outs,
      ins_valid => buffer142_outs_valid,
      ins_ready => buffer142_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork39_outs_0,
      outs(1) => fork39_outs_1,
      outs(2) => fork39_outs_2,
      outs_valid(0) => fork39_outs_0_valid,
      outs_valid(1) => fork39_outs_1_valid,
      outs_valid(2) => fork39_outs_2_valid,
      outs_ready(0) => fork39_outs_0_ready,
      outs_ready(1) => fork39_outs_1_ready,
      outs_ready(2) => fork39_outs_2_ready
    );

  extsi51 : entity work.extsi(arch) generic map(5, 7)
    port map(
      ins => fork39_outs_0,
      ins_valid => fork39_outs_0_valid,
      ins_ready => fork39_outs_0_ready,
      clk => clk,
      rst => rst,
      outs => extsi51_outs,
      outs_valid => extsi51_outs_valid,
      outs_ready => extsi51_outs_ready
    );

  extsi52 : entity work.extsi(arch) generic map(5, 7)
    port map(
      ins => buffer101_outs,
      ins_valid => buffer101_outs_valid,
      ins_ready => buffer101_outs_ready,
      clk => clk,
      rst => rst,
      outs => extsi52_outs,
      outs_valid => extsi52_outs_valid,
      outs_ready => extsi52_outs_ready
    );

  buffer101 : entity work.tfifo(arch) generic map(1, 5)
    port map(
      ins => fork39_outs_1,
      ins_valid => fork39_outs_1_valid,
      ins_ready => fork39_outs_1_ready,
      clk => clk,
      rst => rst,
      outs => buffer101_outs,
      outs_valid => buffer101_outs_valid,
      outs_ready => buffer101_outs_ready
    );

  mux15 : entity work.mux(arch) generic map(2, 32, 1)
    port map(
      index => fork43_outs_2,
      index_valid => fork43_outs_2_valid,
      index_ready => fork43_outs_2_ready,
      ins(0) => buffer130_outs,
      ins(1) => cond_br28_trueOut,
      ins_valid(0) => buffer130_outs_valid,
      ins_valid(1) => cond_br28_trueOut_valid,
      ins_ready(0) => buffer130_outs_ready,
      ins_ready(1) => cond_br28_trueOut_ready,
      clk => clk,
      rst => rst,
      outs => mux15_outs,
      outs_valid => mux15_outs_valid,
      outs_ready => mux15_outs_ready
    );

  buffer145 : entity work.tehb(arch) generic map(32)
    port map(
      ins => mux15_outs,
      ins_valid => mux15_outs_valid,
      ins_ready => mux15_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer145_outs,
      outs_valid => buffer145_outs_valid,
      outs_ready => buffer145_outs_ready
    );

  fork40 : entity work.handshake_fork(arch) generic map(2, 32)
    port map(
      ins => buffer145_outs,
      ins_valid => buffer145_outs_valid,
      ins_ready => buffer145_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork40_outs_0,
      outs(1) => fork40_outs_1,
      outs_valid(0) => fork40_outs_0_valid,
      outs_valid(1) => fork40_outs_1_valid,
      outs_ready(0) => fork40_outs_0_ready,
      outs_ready(1) => fork40_outs_1_ready
    );

  mux16 : entity work.mux(arch) generic map(2, 5, 1)
    port map(
      index => fork43_outs_0,
      index_valid => fork43_outs_0_valid,
      index_ready => fork43_outs_0_ready,
      ins(0) => buffer123_outs,
      ins(1) => cond_br29_trueOut,
      ins_valid(0) => buffer123_outs_valid,
      ins_valid(1) => cond_br29_trueOut_valid,
      ins_ready(0) => buffer123_outs_ready,
      ins_ready(1) => cond_br29_trueOut_ready,
      clk => clk,
      rst => rst,
      outs => mux16_outs,
      outs_valid => mux16_outs_valid,
      outs_ready => mux16_outs_ready
    );

  buffer147 : entity work.oehb(arch) generic map(5)
    port map(
      ins => mux16_outs,
      ins_valid => mux16_outs_valid,
      ins_ready => mux16_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer147_outs,
      outs_valid => buffer147_outs_valid,
      outs_ready => buffer147_outs_ready
    );

  buffer161 : entity work.tehb(arch) generic map(5)
    port map(
      ins => buffer147_outs,
      ins_valid => buffer147_outs_valid,
      ins_ready => buffer147_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer161_outs,
      outs_valid => buffer161_outs_valid,
      outs_ready => buffer161_outs_ready
    );

  fork41 : entity work.handshake_fork(arch) generic map(2, 5)
    port map(
      ins => buffer161_outs,
      ins_valid => buffer161_outs_valid,
      ins_ready => buffer161_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork41_outs_0,
      outs(1) => fork41_outs_1,
      outs_valid(0) => fork41_outs_0_valid,
      outs_valid(1) => fork41_outs_1_valid,
      outs_ready(0) => fork41_outs_0_ready,
      outs_ready(1) => fork41_outs_1_ready
    );

  extsi53 : entity work.extsi(arch) generic map(5, 32)
    port map(
      ins => fork41_outs_1,
      ins_valid => fork41_outs_1_valid,
      ins_ready => fork41_outs_1_ready,
      clk => clk,
      rst => rst,
      outs => extsi53_outs,
      outs_valid => extsi53_outs_valid,
      outs_ready => extsi53_outs_ready
    );

  fork42 : entity work.handshake_fork(arch) generic map(4, 32)
    port map(
      ins => extsi53_outs,
      ins_valid => extsi53_outs_valid,
      ins_ready => extsi53_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork42_outs_0,
      outs(1) => fork42_outs_1,
      outs(2) => fork42_outs_2,
      outs(3) => fork42_outs_3,
      outs_valid(0) => fork42_outs_0_valid,
      outs_valid(1) => fork42_outs_1_valid,
      outs_valid(2) => fork42_outs_2_valid,
      outs_valid(3) => fork42_outs_3_valid,
      outs_ready(0) => fork42_outs_0_ready,
      outs_ready(1) => fork42_outs_1_ready,
      outs_ready(2) => fork42_outs_2_ready,
      outs_ready(3) => fork42_outs_3_ready
    );

  control_merge6 : entity work.control_merge_dataless(arch) generic map(2, 1)
    port map(
      ins_valid(0) => fork35_outs_1_valid,
      ins_valid(1) => cond_br30_trueOut_valid,
      ins_ready(0) => fork35_outs_1_ready,
      ins_ready(1) => cond_br30_trueOut_ready,
      clk => clk,
      rst => rst,
      outs_valid => control_merge6_outs_valid,
      outs_ready => control_merge6_outs_ready,
      index => control_merge6_index,
      index_valid => control_merge6_index_valid,
      index_ready => control_merge6_index_ready
    );

  fork43 : entity work.handshake_fork(arch) generic map(3, 1)
    port map(
      ins => control_merge6_index,
      ins_valid => control_merge6_index_valid,
      ins_ready => control_merge6_index_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork43_outs_0,
      outs(1) => fork43_outs_1,
      outs(2) => fork43_outs_2,
      outs_valid(0) => fork43_outs_0_valid,
      outs_valid(1) => fork43_outs_1_valid,
      outs_valid(2) => fork43_outs_2_valid,
      outs_ready(0) => fork43_outs_0_ready,
      outs_ready(1) => fork43_outs_1_ready,
      outs_ready(2) => fork43_outs_2_ready
    );

  fork44 : entity work.fork_dataless(arch) generic map(3)
    port map(
      ins_valid => control_merge6_outs_valid,
      ins_ready => control_merge6_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid(0) => fork44_outs_0_valid,
      outs_valid(1) => fork44_outs_1_valid,
      outs_valid(2) => fork44_outs_2_valid,
      outs_ready(0) => fork44_outs_0_ready,
      outs_ready(1) => fork44_outs_1_ready,
      outs_ready(2) => fork44_outs_2_ready
    );

  constant45 : entity work.handshake_constant_1(arch) generic map(2)
    port map(
      ctrl_valid => fork44_outs_1_valid,
      ctrl_ready => fork44_outs_1_ready,
      clk => clk,
      rst => rst,
      outs => constant45_outs,
      outs_valid => constant45_outs_valid,
      outs_ready => constant45_outs_ready
    );

  extsi17 : entity work.extsi(arch) generic map(2, 32)
    port map(
      ins => constant45_outs,
      ins_valid => constant45_outs_valid,
      ins_ready => constant45_outs_ready,
      clk => clk,
      rst => rst,
      outs => extsi17_outs,
      outs_valid => extsi17_outs_valid,
      outs_ready => extsi17_outs_ready
    );

  constant46 : entity work.handshake_constant_0(arch) generic map(1)
    port map(
      ctrl_valid => fork44_outs_0_valid,
      ctrl_ready => fork44_outs_0_ready,
      clk => clk,
      rst => rst,
      outs => constant46_outs,
      outs_valid => constant46_outs_valid,
      outs_ready => constant46_outs_ready
    );

  source9 : entity work.source(arch)
    port map(
      clk => clk,
      rst => rst,
      outs_valid => source9_outs_valid,
      outs_ready => source9_outs_ready
    );

  constant47 : entity work.handshake_constant_1(arch) generic map(2)
    port map(
      ctrl_valid => source9_outs_valid,
      ctrl_ready => source9_outs_ready,
      clk => clk,
      rst => rst,
      outs => constant47_outs,
      outs_valid => constant47_outs_valid,
      outs_ready => constant47_outs_ready
    );

  extsi19 : entity work.extsi(arch) generic map(2, 32)
    port map(
      ins => constant47_outs,
      ins_valid => constant47_outs_valid,
      ins_ready => constant47_outs_ready,
      clk => clk,
      rst => rst,
      outs => extsi19_outs,
      outs_valid => extsi19_outs_valid,
      outs_ready => extsi19_outs_ready
    );

  fork45 : entity work.handshake_fork(arch) generic map(2, 32)
    port map(
      ins => extsi19_outs,
      ins_valid => extsi19_outs_valid,
      ins_ready => extsi19_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork45_outs_0,
      outs(1) => fork45_outs_1,
      outs_valid(0) => fork45_outs_0_valid,
      outs_valid(1) => fork45_outs_1_valid,
      outs_ready(0) => fork45_outs_0_ready,
      outs_ready(1) => fork45_outs_1_ready
    );

  source10 : entity work.source(arch)
    port map(
      clk => clk,
      rst => rst,
      outs_valid => source10_outs_valid,
      outs_ready => source10_outs_ready
    );

  constant48 : entity work.handshake_constant_2(arch) generic map(3)
    port map(
      ctrl_valid => source10_outs_valid,
      ctrl_ready => source10_outs_ready,
      clk => clk,
      rst => rst,
      outs => constant48_outs,
      outs_valid => constant48_outs_valid,
      outs_ready => constant48_outs_ready
    );

  extsi20 : entity work.extsi(arch) generic map(3, 32)
    port map(
      ins => constant48_outs,
      ins_valid => constant48_outs_valid,
      ins_ready => constant48_outs_ready,
      clk => clk,
      rst => rst,
      outs => extsi20_outs,
      outs_valid => extsi20_outs_valid,
      outs_ready => extsi20_outs_ready
    );

  fork46 : entity work.handshake_fork(arch) generic map(2, 32)
    port map(
      ins => extsi20_outs,
      ins_valid => extsi20_outs_valid,
      ins_ready => extsi20_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork46_outs_0,
      outs(1) => fork46_outs_1,
      outs_valid(0) => fork46_outs_0_valid,
      outs_valid(1) => fork46_outs_1_valid,
      outs_ready(0) => fork46_outs_0_ready,
      outs_ready(1) => fork46_outs_1_ready
    );

  shli10 : entity work.shli(arch) generic map(32)
    port map(
      lhs => fork42_outs_0,
      lhs_valid => fork42_outs_0_valid,
      lhs_ready => fork42_outs_0_ready,
      rhs => fork45_outs_0,
      rhs_valid => fork45_outs_0_valid,
      rhs_ready => fork45_outs_0_ready,
      clk => clk,
      rst => rst,
      result => shli10_result,
      result_valid => shli10_result_valid,
      result_ready => shli10_result_ready
    );

  buffer163 : entity work.oehb(arch) generic map(32)
    port map(
      ins => shli10_result,
      ins_valid => shli10_result_valid,
      ins_ready => shli10_result_ready,
      clk => clk,
      rst => rst,
      outs => buffer163_outs,
      outs_valid => buffer163_outs_valid,
      outs_ready => buffer163_outs_ready
    );

  trunci11 : entity work.trunci(arch) generic map(32, 7)
    port map(
      ins => buffer163_outs,
      ins_valid => buffer163_outs_valid,
      ins_ready => buffer163_outs_ready,
      clk => clk,
      rst => rst,
      outs => trunci11_outs,
      outs_valid => trunci11_outs_valid,
      outs_ready => trunci11_outs_ready
    );

  shli11 : entity work.shli(arch) generic map(32)
    port map(
      lhs => fork42_outs_1,
      lhs_valid => fork42_outs_1_valid,
      lhs_ready => fork42_outs_1_ready,
      rhs => fork46_outs_0,
      rhs_valid => fork46_outs_0_valid,
      rhs_ready => fork46_outs_0_ready,
      clk => clk,
      rst => rst,
      result => shli11_result,
      result_valid => shli11_result_valid,
      result_ready => shli11_result_ready
    );

  buffer165 : entity work.oehb(arch) generic map(32)
    port map(
      ins => shli11_result,
      ins_valid => shli11_result_valid,
      ins_ready => shli11_result_ready,
      clk => clk,
      rst => rst,
      outs => buffer165_outs,
      outs_valid => buffer165_outs_valid,
      outs_ready => buffer165_outs_ready
    );

  trunci12 : entity work.trunci(arch) generic map(32, 7)
    port map(
      ins => buffer165_outs,
      ins_valid => buffer165_outs_valid,
      ins_ready => buffer165_outs_ready,
      clk => clk,
      rst => rst,
      outs => trunci12_outs,
      outs_valid => trunci12_outs_valid,
      outs_ready => trunci12_outs_ready
    );

  addi24 : entity work.addi(arch) generic map(7)
    port map(
      lhs => trunci11_outs,
      lhs_valid => trunci11_outs_valid,
      lhs_ready => trunci11_outs_ready,
      rhs => trunci12_outs,
      rhs_valid => trunci12_outs_valid,
      rhs_ready => trunci12_outs_ready,
      clk => clk,
      rst => rst,
      result => addi24_result,
      result_valid => addi24_result_valid,
      result_ready => addi24_result_ready
    );

  buffer168 : entity work.oehb(arch) generic map(7)
    port map(
      ins => addi24_result,
      ins_valid => addi24_result_valid,
      ins_ready => addi24_result_ready,
      clk => clk,
      rst => rst,
      outs => buffer168_outs,
      outs_valid => buffer168_outs_valid,
      outs_ready => buffer168_outs_ready
    );

  addi7 : entity work.addi(arch) generic map(7)
    port map(
      lhs => extsi51_outs,
      lhs_valid => extsi51_outs_valid,
      lhs_ready => extsi51_outs_ready,
      rhs => buffer168_outs,
      rhs_valid => buffer168_outs_valid,
      rhs_ready => buffer168_outs_ready,
      clk => clk,
      rst => rst,
      result => addi7_result,
      result_valid => addi7_result_valid,
      result_ready => addi7_result_ready
    );

  buffer2 : entity work.tfifo_dataless(arch) generic map(1)
    port map(
      ins_valid => unbundle2_outs_0_valid,
      ins_ready => unbundle2_outs_0_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer2_outs_valid,
      outs_ready => buffer2_outs_ready
    );

  load3 : entity work.load(arch) generic map(32, 7)
    port map(
      addrIn => addi7_result,
      addrIn_valid => addi7_result_valid,
      addrIn_ready => addi7_result_ready,
      dataFromMem => mem_controller3_ldData_0,
      dataFromMem_valid => mem_controller3_ldData_0_valid,
      dataFromMem_ready => mem_controller3_ldData_0_ready,
      clk => clk,
      rst => rst,
      addrOut => load3_addrOut,
      addrOut_valid => load3_addrOut_valid,
      addrOut_ready => load3_addrOut_ready,
      dataOut => load3_dataOut,
      dataOut_valid => load3_dataOut_valid,
      dataOut_ready => load3_dataOut_ready
    );

  fork47 : entity work.handshake_fork(arch) generic map(2, 32)
    port map(
      ins => load3_dataOut,
      ins_valid => load3_dataOut_valid,
      ins_ready => load3_dataOut_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork47_outs_0,
      outs(1) => fork47_outs_1,
      outs_valid(0) => fork47_outs_0_valid,
      outs_valid(1) => fork47_outs_1_valid,
      outs_ready(0) => fork47_outs_0_ready,
      outs_ready(1) => fork47_outs_1_ready
    );

  muli2 : entity work.muli(arch) generic map(32)
    port map(
      lhs => fork47_outs_1,
      lhs_valid => fork47_outs_1_valid,
      lhs_ready => fork47_outs_1_ready,
      rhs => buffer110_outs,
      rhs_valid => buffer110_outs_valid,
      rhs_ready => buffer110_outs_ready,
      clk => clk,
      rst => rst,
      result => muli2_result,
      result_valid => muli2_result_valid,
      result_ready => muli2_result_ready
    );

  buffer110 : entity work.tfifo(arch) generic map(1, 32)
    port map(
      ins => fork40_outs_1,
      ins_valid => fork40_outs_1_valid,
      ins_ready => fork40_outs_1_ready,
      clk => clk,
      rst => rst,
      outs => buffer110_outs,
      outs_valid => buffer110_outs_valid,
      outs_ready => buffer110_outs_ready
    );

  shli12 : entity work.shli(arch) generic map(32)
    port map(
      lhs => buffer112_outs,
      lhs_valid => buffer112_outs_valid,
      lhs_ready => buffer112_outs_ready,
      rhs => buffer111_outs,
      rhs_valid => buffer111_outs_valid,
      rhs_ready => buffer111_outs_ready,
      clk => clk,
      rst => rst,
      result => shli12_result,
      result_valid => shli12_result_valid,
      result_ready => shli12_result_ready
    );

  buffer111 : entity work.tfifo(arch) generic map(1, 32)
    port map(
      ins => fork45_outs_1,
      ins_valid => fork45_outs_1_valid,
      ins_ready => fork45_outs_1_ready,
      clk => clk,
      rst => rst,
      outs => buffer111_outs,
      outs_valid => buffer111_outs_valid,
      outs_ready => buffer111_outs_ready
    );

  buffer112 : entity work.tfifo(arch) generic map(1, 32)
    port map(
      ins => fork42_outs_2,
      ins_valid => fork42_outs_2_valid,
      ins_ready => fork42_outs_2_ready,
      clk => clk,
      rst => rst,
      outs => buffer112_outs,
      outs_valid => buffer112_outs_valid,
      outs_ready => buffer112_outs_ready
    );

  buffer171 : entity work.oehb(arch) generic map(32)
    port map(
      ins => shli12_result,
      ins_valid => shli12_result_valid,
      ins_ready => shli12_result_ready,
      clk => clk,
      rst => rst,
      outs => buffer171_outs,
      outs_valid => buffer171_outs_valid,
      outs_ready => buffer171_outs_ready
    );

  trunci13 : entity work.trunci(arch) generic map(32, 7)
    port map(
      ins => buffer171_outs,
      ins_valid => buffer171_outs_valid,
      ins_ready => buffer171_outs_ready,
      clk => clk,
      rst => rst,
      outs => trunci13_outs,
      outs_valid => trunci13_outs_valid,
      outs_ready => trunci13_outs_ready
    );

  shli13 : entity work.shli(arch) generic map(32)
    port map(
      lhs => fork42_outs_3,
      lhs_valid => fork42_outs_3_valid,
      lhs_ready => fork42_outs_3_ready,
      rhs => buffer113_outs,
      rhs_valid => buffer113_outs_valid,
      rhs_ready => buffer113_outs_ready,
      clk => clk,
      rst => rst,
      result => shli13_result,
      result_valid => shli13_result_valid,
      result_ready => shli13_result_ready
    );

  buffer113 : entity work.tfifo(arch) generic map(1, 32)
    port map(
      ins => fork46_outs_1,
      ins_valid => fork46_outs_1_valid,
      ins_ready => fork46_outs_1_ready,
      clk => clk,
      rst => rst,
      outs => buffer113_outs,
      outs_valid => buffer113_outs_valid,
      outs_ready => buffer113_outs_ready
    );

  buffer172 : entity work.oehb(arch) generic map(32)
    port map(
      ins => shli13_result,
      ins_valid => shli13_result_valid,
      ins_ready => shli13_result_ready,
      clk => clk,
      rst => rst,
      outs => buffer172_outs,
      outs_valid => buffer172_outs_valid,
      outs_ready => buffer172_outs_ready
    );

  trunci14 : entity work.trunci(arch) generic map(32, 7)
    port map(
      ins => buffer172_outs,
      ins_valid => buffer172_outs_valid,
      ins_ready => buffer172_outs_ready,
      clk => clk,
      rst => rst,
      outs => trunci14_outs,
      outs_valid => trunci14_outs_valid,
      outs_ready => trunci14_outs_ready
    );

  addi25 : entity work.addi(arch) generic map(7)
    port map(
      lhs => trunci13_outs,
      lhs_valid => trunci13_outs_valid,
      lhs_ready => trunci13_outs_ready,
      rhs => trunci14_outs,
      rhs_valid => trunci14_outs_valid,
      rhs_ready => trunci14_outs_ready,
      clk => clk,
      rst => rst,
      result => addi25_result,
      result_valid => addi25_result_valid,
      result_ready => addi25_result_ready
    );

  buffer173 : entity work.oehb(arch) generic map(7)
    port map(
      ins => addi25_result,
      ins_valid => addi25_result_valid,
      ins_ready => addi25_result_ready,
      clk => clk,
      rst => rst,
      outs => buffer173_outs,
      outs_valid => buffer173_outs_valid,
      outs_ready => buffer173_outs_ready
    );

  addi8 : entity work.addi(arch) generic map(7)
    port map(
      lhs => extsi52_outs,
      lhs_valid => extsi52_outs_valid,
      lhs_ready => extsi52_outs_ready,
      rhs => buffer173_outs,
      rhs_valid => buffer173_outs_valid,
      rhs_ready => buffer173_outs_ready,
      clk => clk,
      rst => rst,
      result => addi8_result,
      result_valid => addi8_result_valid,
      result_ready => addi8_result_ready
    );

  buffer3 : entity work.tfifo_dataless(arch) generic map(1)
    port map(
      ins_valid => store2_doneOut_valid,
      ins_ready => store2_doneOut_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer3_outs_valid,
      outs_ready => buffer3_outs_ready
    );

  buffer175 : entity work.oehb(arch) generic map(7)
    port map(
      ins => addi8_result,
      ins_valid => addi8_result_valid,
      ins_ready => addi8_result_ready,
      clk => clk,
      rst => rst,
      outs => buffer175_outs,
      outs_valid => buffer175_outs_valid,
      outs_ready => buffer175_outs_ready
    );

  store2 : entity work.store(arch) generic map(32, 7)
    port map(
      addrIn => buffer175_outs,
      addrIn_valid => buffer175_outs_valid,
      addrIn_ready => buffer175_outs_ready,
      dataIn => muli2_result,
      dataIn_valid => muli2_result_valid,
      dataIn_ready => muli2_result_ready,
      doneFromMem_valid => mem_controller3_stDone_0_valid,
      doneFromMem_ready => mem_controller3_stDone_0_ready,
      clk => clk,
      rst => rst,
      addrOut => store2_addrOut,
      addrOut_valid => store2_addrOut_valid,
      addrOut_ready => store2_addrOut_ready,
      dataToMem => store2_dataToMem,
      dataToMem_valid => store2_dataToMem_valid,
      dataToMem_ready => store2_dataToMem_ready,
      doneOut_valid => store2_doneOut_valid,
      doneOut_ready => store2_doneOut_ready
    );

  extsi29 : entity work.extsi(arch) generic map(1, 5)
    port map(
      ins => constant46_outs,
      ins_valid => constant46_outs_valid,
      ins_ready => constant46_outs_ready,
      clk => clk,
      rst => rst,
      outs => extsi29_outs,
      outs_valid => extsi29_outs_valid,
      outs_ready => extsi29_outs_ready
    );

  cond_br89 : entity work.cond_br_dataless(arch)
    port map(
      condition => buffer118_outs,
      condition_valid => buffer118_outs_valid,
      condition_ready => buffer118_outs_ready,
      data_valid => fork50_outs_1_valid,
      data_ready => fork50_outs_1_ready,
      clk => clk,
      rst => rst,
      trueOut_valid => cond_br89_trueOut_valid,
      trueOut_ready => cond_br89_trueOut_ready,
      falseOut_valid => cond_br89_falseOut_valid,
      falseOut_ready => cond_br89_falseOut_ready
    );

  buffer118 : entity work.tfifo(arch) generic map(1, 1)
    port map(
      ins => fork65_outs_8,
      ins_valid => fork65_outs_8_valid,
      ins_ready => fork65_outs_8_ready,
      clk => clk,
      rst => rst,
      outs => buffer118_outs,
      outs_valid => buffer118_outs_valid,
      outs_ready => buffer118_outs_ready
    );

  sink10 : entity work.sink_dataless(arch)
    port map(
      ins_valid => cond_br89_falseOut_valid,
      ins_ready => cond_br89_falseOut_ready,
      clk => clk,
      rst => rst
    );

  cond_br90 : entity work.cond_br_dataless(arch)
    port map(
      condition => buffer119_outs,
      condition_valid => buffer119_outs_valid,
      condition_ready => buffer119_outs_ready,
      data_valid => fork52_outs_1_valid,
      data_ready => fork52_outs_1_ready,
      clk => clk,
      rst => rst,
      trueOut_valid => cond_br90_trueOut_valid,
      trueOut_ready => cond_br90_trueOut_ready,
      falseOut_valid => cond_br90_falseOut_valid,
      falseOut_ready => cond_br90_falseOut_ready
    );

  buffer119 : entity work.tfifo(arch) generic map(4, 1)
    port map(
      ins => fork65_outs_7,
      ins_valid => fork65_outs_7_valid,
      ins_ready => fork65_outs_7_ready,
      clk => clk,
      rst => rst,
      outs => buffer119_outs,
      outs_valid => buffer119_outs_valid,
      outs_ready => buffer119_outs_ready
    );

  sink11 : entity work.sink_dataless(arch)
    port map(
      ins_valid => cond_br90_falseOut_valid,
      ins_ready => cond_br90_falseOut_ready,
      clk => clk,
      rst => rst
    );

  cond_br91 : entity work.cond_br_dataless(arch)
    port map(
      condition => buffer120_outs,
      condition_valid => buffer120_outs_valid,
      condition_ready => buffer120_outs_ready,
      data_valid => fork49_outs_2_valid,
      data_ready => fork49_outs_2_ready,
      clk => clk,
      rst => rst,
      trueOut_valid => cond_br91_trueOut_valid,
      trueOut_ready => cond_br91_trueOut_ready,
      falseOut_valid => cond_br91_falseOut_valid,
      falseOut_ready => cond_br91_falseOut_ready
    );

  buffer120 : entity work.tfifo(arch) generic map(3, 1)
    port map(
      ins => fork65_outs_6,
      ins_valid => fork65_outs_6_valid,
      ins_ready => fork65_outs_6_ready,
      clk => clk,
      rst => rst,
      outs => buffer120_outs,
      outs_valid => buffer120_outs_valid,
      outs_ready => buffer120_outs_ready
    );

  sink12 : entity work.sink_dataless(arch)
    port map(
      ins_valid => cond_br91_falseOut_valid,
      ins_ready => cond_br91_falseOut_ready,
      clk => clk,
      rst => rst
    );

  cond_br92 : entity work.cond_br_dataless(arch)
    port map(
      condition => fork65_outs_5,
      condition_valid => fork65_outs_5_valid,
      condition_ready => fork65_outs_5_ready,
      data_valid => fork51_outs_1_valid,
      data_ready => fork51_outs_1_ready,
      clk => clk,
      rst => rst,
      trueOut_valid => cond_br92_trueOut_valid,
      trueOut_ready => cond_br92_trueOut_ready,
      falseOut_valid => cond_br92_falseOut_valid,
      falseOut_ready => cond_br92_falseOut_ready
    );

  sink13 : entity work.sink_dataless(arch)
    port map(
      ins_valid => cond_br92_falseOut_valid,
      ins_ready => cond_br92_falseOut_ready,
      clk => clk,
      rst => rst
    );

  buffer209 : entity work.oehb_dataless(arch)
    port map(
      ins_valid => buffer4_outs_valid,
      ins_ready => buffer4_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer209_outs_valid,
      outs_ready => buffer209_outs_ready
    );

  cond_br93 : entity work.cond_br_dataless(arch)
    port map(
      condition => buffer122_outs,
      condition_valid => buffer122_outs_valid,
      condition_ready => buffer122_outs_ready,
      data_valid => buffer209_outs_valid,
      data_ready => buffer209_outs_ready,
      clk => clk,
      rst => rst,
      trueOut_valid => cond_br93_trueOut_valid,
      trueOut_ready => cond_br93_trueOut_ready,
      falseOut_valid => cond_br93_falseOut_valid,
      falseOut_ready => cond_br93_falseOut_ready
    );

  buffer122 : entity work.tfifo(arch) generic map(4, 1)
    port map(
      ins => fork65_outs_4,
      ins_valid => fork65_outs_4_valid,
      ins_ready => fork65_outs_4_ready,
      clk => clk,
      rst => rst,
      outs => buffer122_outs,
      outs_valid => buffer122_outs_valid,
      outs_ready => buffer122_outs_ready
    );

  init26 : entity work.tehb_init(arch) generic map(1, 0)
    port map(
      ins => fork65_outs_3,
      ins_valid => fork65_outs_3_valid,
      ins_ready => fork65_outs_3_ready,
      clk => clk,
      rst => rst,
      outs => init26_outs,
      outs_valid => init26_outs_valid,
      outs_ready => init26_outs_ready
    );

  fork48 : entity work.handshake_fork(arch) generic map(5, 1)
    port map(
      ins => init26_outs,
      ins_valid => init26_outs_valid,
      ins_ready => init26_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork48_outs_0,
      outs(1) => fork48_outs_1,
      outs(2) => fork48_outs_2,
      outs(3) => fork48_outs_3,
      outs(4) => fork48_outs_4,
      outs_valid(0) => fork48_outs_0_valid,
      outs_valid(1) => fork48_outs_1_valid,
      outs_valid(2) => fork48_outs_2_valid,
      outs_valid(3) => fork48_outs_3_valid,
      outs_valid(4) => fork48_outs_4_valid,
      outs_ready(0) => fork48_outs_0_ready,
      outs_ready(1) => fork48_outs_1_ready,
      outs_ready(2) => fork48_outs_2_ready,
      outs_ready(3) => fork48_outs_3_ready,
      outs_ready(4) => fork48_outs_4_ready
    );

  mux47 : entity work.mux_dataless(arch) generic map(2, 1)
    port map(
      index => buffer124_outs,
      index_valid => buffer124_outs_valid,
      index_ready => buffer124_outs_ready,
      ins_valid(0) => buffer3_outs_valid,
      ins_valid(1) => cond_br91_trueOut_valid,
      ins_ready(0) => buffer3_outs_ready,
      ins_ready(1) => cond_br91_trueOut_ready,
      clk => clk,
      rst => rst,
      outs_valid => mux47_outs_valid,
      outs_ready => mux47_outs_ready
    );

  buffer124 : entity work.tfifo(arch) generic map(3, 1)
    port map(
      ins => fork48_outs_4,
      ins_valid => fork48_outs_4_valid,
      ins_ready => fork48_outs_4_ready,
      clk => clk,
      rst => rst,
      outs => buffer124_outs,
      outs_valid => buffer124_outs_valid,
      outs_ready => buffer124_outs_ready
    );

  buffer178 : entity work.oehb_dataless(arch)
    port map(
      ins_valid => mux47_outs_valid,
      ins_ready => mux47_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer178_outs_valid,
      outs_ready => buffer178_outs_ready
    );

  buffer179 : entity work.tehb_dataless(arch)
    port map(
      ins_valid => buffer178_outs_valid,
      ins_ready => buffer178_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer179_outs_valid,
      outs_ready => buffer179_outs_ready
    );

  fork49 : entity work.fork_dataless(arch) generic map(3)
    port map(
      ins_valid => buffer179_outs_valid,
      ins_ready => buffer179_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid(0) => fork49_outs_0_valid,
      outs_valid(1) => fork49_outs_1_valid,
      outs_valid(2) => fork49_outs_2_valid,
      outs_ready(0) => fork49_outs_0_ready,
      outs_ready(1) => fork49_outs_1_ready,
      outs_ready(2) => fork49_outs_2_ready
    );

  mux48 : entity work.mux_dataless(arch) generic map(2, 1)
    port map(
      index => buffer125_outs,
      index_valid => buffer125_outs_valid,
      index_ready => buffer125_outs_ready,
      ins_valid(0) => fork37_outs_1_valid,
      ins_valid(1) => cond_br89_trueOut_valid,
      ins_ready(0) => fork37_outs_1_ready,
      ins_ready(1) => cond_br89_trueOut_ready,
      clk => clk,
      rst => rst,
      outs_valid => mux48_outs_valid,
      outs_ready => mux48_outs_ready
    );

  buffer125 : entity work.tfifo(arch) generic map(1, 1)
    port map(
      ins => fork48_outs_3,
      ins_valid => fork48_outs_3_valid,
      ins_ready => fork48_outs_3_ready,
      clk => clk,
      rst => rst,
      outs => buffer125_outs,
      outs_valid => buffer125_outs_valid,
      outs_ready => buffer125_outs_ready
    );

  buffer180 : entity work.oehb_dataless(arch)
    port map(
      ins_valid => mux48_outs_valid,
      ins_ready => mux48_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer180_outs_valid,
      outs_ready => buffer180_outs_ready
    );

  buffer181 : entity work.tehb_dataless(arch)
    port map(
      ins_valid => buffer180_outs_valid,
      ins_ready => buffer180_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer181_outs_valid,
      outs_ready => buffer181_outs_ready
    );

  fork50 : entity work.fork_dataless(arch) generic map(2)
    port map(
      ins_valid => buffer181_outs_valid,
      ins_ready => buffer181_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid(0) => fork50_outs_0_valid,
      outs_valid(1) => fork50_outs_1_valid,
      outs_ready(0) => fork50_outs_0_ready,
      outs_ready(1) => fork50_outs_1_ready
    );

  mux49 : entity work.mux_dataless(arch) generic map(2, 1)
    port map(
      index => buffer126_outs,
      index_valid => buffer126_outs_valid,
      index_ready => buffer126_outs_ready,
      ins_valid(0) => fork38_outs_1_valid,
      ins_valid(1) => cond_br92_trueOut_valid,
      ins_ready(0) => fork38_outs_1_ready,
      ins_ready(1) => cond_br92_trueOut_ready,
      clk => clk,
      rst => rst,
      outs_valid => mux49_outs_valid,
      outs_ready => mux49_outs_ready
    );

  buffer126 : entity work.tfifo(arch) generic map(1, 1)
    port map(
      ins => fork48_outs_2,
      ins_valid => fork48_outs_2_valid,
      ins_ready => fork48_outs_2_ready,
      clk => clk,
      rst => rst,
      outs => buffer126_outs,
      outs_valid => buffer126_outs_valid,
      outs_ready => buffer126_outs_ready
    );

  buffer182 : entity work.oehb_dataless(arch)
    port map(
      ins_valid => mux49_outs_valid,
      ins_ready => mux49_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer182_outs_valid,
      outs_ready => buffer182_outs_ready
    );

  buffer183 : entity work.tehb_dataless(arch)
    port map(
      ins_valid => buffer182_outs_valid,
      ins_ready => buffer182_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer183_outs_valid,
      outs_ready => buffer183_outs_ready
    );

  fork51 : entity work.fork_dataless(arch) generic map(2)
    port map(
      ins_valid => buffer183_outs_valid,
      ins_ready => buffer183_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid(0) => fork51_outs_0_valid,
      outs_valid(1) => fork51_outs_1_valid,
      outs_ready(0) => fork51_outs_0_ready,
      outs_ready(1) => fork51_outs_1_ready
    );

  mux51 : entity work.mux_dataless(arch) generic map(2, 1)
    port map(
      index => buffer127_outs,
      index_valid => buffer127_outs_valid,
      index_ready => buffer127_outs_ready,
      ins_valid(0) => buffer2_outs_valid,
      ins_valid(1) => cond_br90_trueOut_valid,
      ins_ready(0) => buffer2_outs_ready,
      ins_ready(1) => cond_br90_trueOut_ready,
      clk => clk,
      rst => rst,
      outs_valid => mux51_outs_valid,
      outs_ready => mux51_outs_ready
    );

  buffer127 : entity work.tfifo(arch) generic map(3, 1)
    port map(
      ins => fork48_outs_1,
      ins_valid => fork48_outs_1_valid,
      ins_ready => fork48_outs_1_ready,
      clk => clk,
      rst => rst,
      outs => buffer127_outs,
      outs_valid => buffer127_outs_valid,
      outs_ready => buffer127_outs_ready
    );

  buffer185 : entity work.oehb_dataless(arch)
    port map(
      ins_valid => mux51_outs_valid,
      ins_ready => mux51_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer185_outs_valid,
      outs_ready => buffer185_outs_ready
    );

  buffer186 : entity work.tehb_dataless(arch)
    port map(
      ins_valid => buffer185_outs_valid,
      ins_ready => buffer185_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer186_outs_valid,
      outs_ready => buffer186_outs_ready
    );

  fork52 : entity work.fork_dataless(arch) generic map(2)
    port map(
      ins_valid => buffer186_outs_valid,
      ins_ready => buffer186_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid(0) => fork52_outs_0_valid,
      outs_valid(1) => fork52_outs_1_valid,
      outs_ready(0) => fork52_outs_0_ready,
      outs_ready(1) => fork52_outs_1_ready
    );

  buffer136 : entity work.oehb_dataless(arch)
    port map(
      ins_valid => mux46_outs_valid,
      ins_ready => mux46_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer136_outs_valid,
      outs_ready => buffer136_outs_ready
    );

  buffer140 : entity work.tehb_dataless(arch)
    port map(
      ins_valid => buffer136_outs_valid,
      ins_ready => buffer136_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer140_outs_valid,
      outs_ready => buffer140_outs_ready
    );

  mux52 : entity work.mux_dataless(arch) generic map(2, 1)
    port map(
      index => buffer128_outs,
      index_valid => buffer128_outs_valid,
      index_ready => buffer128_outs_ready,
      ins_valid(0) => buffer140_outs_valid,
      ins_valid(1) => cond_br93_trueOut_valid,
      ins_ready(0) => buffer140_outs_ready,
      ins_ready(1) => cond_br93_trueOut_ready,
      clk => clk,
      rst => rst,
      outs_valid => mux52_outs_valid,
      outs_ready => mux52_outs_ready
    );

  buffer128 : entity work.tfifo(arch) generic map(3, 1)
    port map(
      ins => fork48_outs_0,
      ins_valid => fork48_outs_0_valid,
      ins_ready => fork48_outs_0_ready,
      clk => clk,
      rst => rst,
      outs => buffer128_outs,
      outs_valid => buffer128_outs_valid,
      outs_ready => buffer128_outs_ready
    );

  mux17 : entity work.mux(arch) generic map(2, 5, 1)
    port map(
      index => fork59_outs_2,
      index_valid => fork59_outs_2_valid,
      index_ready => fork59_outs_2_ready,
      ins(0) => extsi29_outs,
      ins(1) => cond_br22_trueOut,
      ins_valid(0) => extsi29_outs_valid,
      ins_valid(1) => cond_br22_trueOut_valid,
      ins_ready(0) => extsi29_outs_ready,
      ins_ready(1) => cond_br22_trueOut_ready,
      clk => clk,
      rst => rst,
      outs => mux17_outs,
      outs_valid => mux17_outs_valid,
      outs_ready => mux17_outs_ready
    );

  buffer188 : entity work.oehb(arch) generic map(5)
    port map(
      ins => mux17_outs,
      ins_valid => mux17_outs_valid,
      ins_ready => mux17_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer188_outs,
      outs_valid => buffer188_outs_valid,
      outs_ready => buffer188_outs_ready
    );

  buffer189 : entity work.tehb(arch) generic map(5)
    port map(
      ins => buffer188_outs,
      ins_valid => buffer188_outs_valid,
      ins_ready => buffer188_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer189_outs,
      outs_valid => buffer189_outs_valid,
      outs_ready => buffer189_outs_ready
    );

  fork53 : entity work.handshake_fork(arch) generic map(2, 5)
    port map(
      ins => buffer189_outs,
      ins_valid => buffer189_outs_valid,
      ins_ready => buffer189_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork53_outs_0,
      outs(1) => fork53_outs_1,
      outs_valid(0) => fork53_outs_0_valid,
      outs_valid(1) => fork53_outs_1_valid,
      outs_ready(0) => fork53_outs_0_ready,
      outs_ready(1) => fork53_outs_1_ready
    );

  extsi54 : entity work.extsi(arch) generic map(5, 6)
    port map(
      ins => fork53_outs_0,
      ins_valid => fork53_outs_0_valid,
      ins_ready => fork53_outs_0_ready,
      clk => clk,
      rst => rst,
      outs => extsi54_outs,
      outs_valid => extsi54_outs_valid,
      outs_ready => extsi54_outs_ready
    );

  extsi55 : entity work.extsi(arch) generic map(5, 32)
    port map(
      ins => fork53_outs_1,
      ins_valid => fork53_outs_1_valid,
      ins_ready => fork53_outs_1_ready,
      clk => clk,
      rst => rst,
      outs => extsi55_outs,
      outs_valid => extsi55_outs_valid,
      outs_ready => extsi55_outs_ready
    );

  fork54 : entity work.handshake_fork(arch) generic map(3, 32)
    port map(
      ins => extsi55_outs,
      ins_valid => extsi55_outs_valid,
      ins_ready => extsi55_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork54_outs_0,
      outs(1) => fork54_outs_1,
      outs(2) => fork54_outs_2,
      outs_valid(0) => fork54_outs_0_valid,
      outs_valid(1) => fork54_outs_1_valid,
      outs_valid(2) => fork54_outs_2_valid,
      outs_ready(0) => fork54_outs_0_ready,
      outs_ready(1) => fork54_outs_1_ready,
      outs_ready(2) => fork54_outs_2_ready
    );

  mux18 : entity work.mux(arch) generic map(2, 32, 1)
    port map(
      index => fork59_outs_3,
      index_valid => fork59_outs_3_valid,
      index_ready => fork59_outs_3_ready,
      ins(0) => fork40_outs_0,
      ins(1) => cond_br23_trueOut,
      ins_valid(0) => fork40_outs_0_valid,
      ins_valid(1) => cond_br23_trueOut_valid,
      ins_ready(0) => fork40_outs_0_ready,
      ins_ready(1) => cond_br23_trueOut_ready,
      clk => clk,
      rst => rst,
      outs => mux18_outs,
      outs_valid => mux18_outs_valid,
      outs_ready => mux18_outs_ready
    );

  mux19 : entity work.mux(arch) generic map(2, 5, 1)
    port map(
      index => fork59_outs_0,
      index_valid => fork59_outs_0_valid,
      index_ready => fork59_outs_0_ready,
      ins(0) => fork41_outs_0,
      ins(1) => cond_br24_trueOut,
      ins_valid(0) => fork41_outs_0_valid,
      ins_valid(1) => cond_br24_trueOut_valid,
      ins_ready(0) => fork41_outs_0_ready,
      ins_ready(1) => cond_br24_trueOut_ready,
      clk => clk,
      rst => rst,
      outs => mux19_outs,
      outs_valid => mux19_outs_valid,
      outs_ready => mux19_outs_ready
    );

  buffer192 : entity work.oehb(arch) generic map(5)
    port map(
      ins => mux19_outs,
      ins_valid => mux19_outs_valid,
      ins_ready => mux19_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer192_outs,
      outs_valid => buffer192_outs_valid,
      outs_ready => buffer192_outs_ready
    );

  buffer193 : entity work.tehb(arch) generic map(5)
    port map(
      ins => buffer192_outs,
      ins_valid => buffer192_outs_valid,
      ins_ready => buffer192_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer193_outs,
      outs_valid => buffer193_outs_valid,
      outs_ready => buffer193_outs_ready
    );

  fork55 : entity work.handshake_fork(arch) generic map(2, 5)
    port map(
      ins => buffer193_outs,
      ins_valid => buffer193_outs_valid,
      ins_ready => buffer193_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork55_outs_0,
      outs(1) => fork55_outs_1,
      outs_valid(0) => fork55_outs_0_valid,
      outs_valid(1) => fork55_outs_1_valid,
      outs_ready(0) => fork55_outs_0_ready,
      outs_ready(1) => fork55_outs_1_ready
    );

  extsi56 : entity work.extsi(arch) generic map(5, 32)
    port map(
      ins => buffer134_outs,
      ins_valid => buffer134_outs_valid,
      ins_ready => buffer134_outs_ready,
      clk => clk,
      rst => rst,
      outs => extsi56_outs,
      outs_valid => extsi56_outs_valid,
      outs_ready => extsi56_outs_ready
    );

  buffer134 : entity work.tfifo(arch) generic map(1, 5)
    port map(
      ins => fork55_outs_1,
      ins_valid => fork55_outs_1_valid,
      ins_ready => fork55_outs_1_ready,
      clk => clk,
      rst => rst,
      outs => buffer134_outs,
      outs_valid => buffer134_outs_valid,
      outs_ready => buffer134_outs_ready
    );

  fork56 : entity work.handshake_fork(arch) generic map(6, 32)
    port map(
      ins => extsi56_outs,
      ins_valid => extsi56_outs_valid,
      ins_ready => extsi56_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork56_outs_0,
      outs(1) => fork56_outs_1,
      outs(2) => fork56_outs_2,
      outs(3) => fork56_outs_3,
      outs(4) => fork56_outs_4,
      outs(5) => fork56_outs_5,
      outs_valid(0) => fork56_outs_0_valid,
      outs_valid(1) => fork56_outs_1_valid,
      outs_valid(2) => fork56_outs_2_valid,
      outs_valid(3) => fork56_outs_3_valid,
      outs_valid(4) => fork56_outs_4_valid,
      outs_valid(5) => fork56_outs_5_valid,
      outs_ready(0) => fork56_outs_0_ready,
      outs_ready(1) => fork56_outs_1_ready,
      outs_ready(2) => fork56_outs_2_ready,
      outs_ready(3) => fork56_outs_3_ready,
      outs_ready(4) => fork56_outs_4_ready,
      outs_ready(5) => fork56_outs_5_ready
    );

  mux20 : entity work.mux(arch) generic map(2, 5, 1)
    port map(
      index => fork59_outs_1,
      index_valid => fork59_outs_1_valid,
      index_ready => fork59_outs_1_ready,
      ins(0) => fork39_outs_2,
      ins(1) => cond_br25_trueOut,
      ins_valid(0) => fork39_outs_2_valid,
      ins_valid(1) => cond_br25_trueOut_valid,
      ins_ready(0) => fork39_outs_2_ready,
      ins_ready(1) => cond_br25_trueOut_ready,
      clk => clk,
      rst => rst,
      outs => mux20_outs,
      outs_valid => mux20_outs_valid,
      outs_ready => mux20_outs_ready
    );

  buffer194 : entity work.oehb(arch) generic map(5)
    port map(
      ins => mux20_outs,
      ins_valid => mux20_outs_valid,
      ins_ready => mux20_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer194_outs,
      outs_valid => buffer194_outs_valid,
      outs_ready => buffer194_outs_ready
    );

  buffer195 : entity work.tehb(arch) generic map(5)
    port map(
      ins => buffer194_outs,
      ins_valid => buffer194_outs_valid,
      ins_ready => buffer194_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer195_outs,
      outs_valid => buffer195_outs_valid,
      outs_ready => buffer195_outs_ready
    );

  fork57 : entity work.handshake_fork(arch) generic map(3, 5)
    port map(
      ins => buffer195_outs,
      ins_valid => buffer195_outs_valid,
      ins_ready => buffer195_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork57_outs_0,
      outs(1) => fork57_outs_1,
      outs(2) => fork57_outs_2,
      outs_valid(0) => fork57_outs_0_valid,
      outs_valid(1) => fork57_outs_1_valid,
      outs_valid(2) => fork57_outs_2_valid,
      outs_ready(0) => fork57_outs_0_ready,
      outs_ready(1) => fork57_outs_1_ready,
      outs_ready(2) => fork57_outs_2_ready
    );

  extsi57 : entity work.extsi(arch) generic map(5, 7)
    port map(
      ins => fork57_outs_0,
      ins_valid => fork57_outs_0_valid,
      ins_ready => fork57_outs_0_ready,
      clk => clk,
      rst => rst,
      outs => extsi57_outs,
      outs_valid => extsi57_outs_valid,
      outs_ready => extsi57_outs_ready
    );

  extsi58 : entity work.extsi(arch) generic map(5, 32)
    port map(
      ins => buffer137_outs,
      ins_valid => buffer137_outs_valid,
      ins_ready => buffer137_outs_ready,
      clk => clk,
      rst => rst,
      outs => extsi58_outs,
      outs_valid => extsi58_outs_valid,
      outs_ready => extsi58_outs_ready
    );

  buffer137 : entity work.tfifo(arch) generic map(1, 5)
    port map(
      ins => fork57_outs_2,
      ins_valid => fork57_outs_2_valid,
      ins_ready => fork57_outs_2_ready,
      clk => clk,
      rst => rst,
      outs => buffer137_outs,
      outs_valid => buffer137_outs_valid,
      outs_ready => buffer137_outs_ready
    );

  fork58 : entity work.handshake_fork(arch) generic map(2, 32)
    port map(
      ins => extsi58_outs,
      ins_valid => extsi58_outs_valid,
      ins_ready => extsi58_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork58_outs_0,
      outs(1) => fork58_outs_1,
      outs_valid(0) => fork58_outs_0_valid,
      outs_valid(1) => fork58_outs_1_valid,
      outs_ready(0) => fork58_outs_0_ready,
      outs_ready(1) => fork58_outs_1_ready
    );

  control_merge7 : entity work.control_merge_dataless(arch) generic map(2, 1)
    port map(
      ins_valid(0) => fork44_outs_2_valid,
      ins_valid(1) => cond_br26_trueOut_valid,
      ins_ready(0) => fork44_outs_2_ready,
      ins_ready(1) => cond_br26_trueOut_ready,
      clk => clk,
      rst => rst,
      outs_valid => control_merge7_outs_valid,
      outs_ready => control_merge7_outs_ready,
      index => control_merge7_index,
      index_valid => control_merge7_index_valid,
      index_ready => control_merge7_index_ready
    );

  fork59 : entity work.handshake_fork(arch) generic map(4, 1)
    port map(
      ins => control_merge7_index,
      ins_valid => control_merge7_index_valid,
      ins_ready => control_merge7_index_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork59_outs_0,
      outs(1) => fork59_outs_1,
      outs(2) => fork59_outs_2,
      outs(3) => fork59_outs_3,
      outs_valid(0) => fork59_outs_0_valid,
      outs_valid(1) => fork59_outs_1_valid,
      outs_valid(2) => fork59_outs_2_valid,
      outs_valid(3) => fork59_outs_3_valid,
      outs_ready(0) => fork59_outs_0_ready,
      outs_ready(1) => fork59_outs_1_ready,
      outs_ready(2) => fork59_outs_2_ready,
      outs_ready(3) => fork59_outs_3_ready
    );

  buffer196 : entity work.oehb_dataless(arch)
    port map(
      ins_valid => control_merge7_outs_valid,
      ins_ready => control_merge7_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer196_outs_valid,
      outs_ready => buffer196_outs_ready
    );

  fork60 : entity work.fork_dataless(arch) generic map(2)
    port map(
      ins_valid => buffer196_outs_valid,
      ins_ready => buffer196_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid(0) => fork60_outs_0_valid,
      outs_valid(1) => fork60_outs_1_valid,
      outs_ready(0) => fork60_outs_0_ready,
      outs_ready(1) => fork60_outs_1_ready
    );

  constant49 : entity work.handshake_constant_1(arch) generic map(2)
    port map(
      ctrl_valid => fork60_outs_0_valid,
      ctrl_ready => fork60_outs_0_ready,
      clk => clk,
      rst => rst,
      outs => constant49_outs,
      outs_valid => constant49_outs_valid,
      outs_ready => constant49_outs_ready
    );

  extsi21 : entity work.extsi(arch) generic map(2, 32)
    port map(
      ins => constant49_outs,
      ins_valid => constant49_outs_valid,
      ins_ready => constant49_outs_ready,
      clk => clk,
      rst => rst,
      outs => extsi21_outs,
      outs_valid => extsi21_outs_valid,
      outs_ready => extsi21_outs_ready
    );

  source11 : entity work.source(arch)
    port map(
      clk => clk,
      rst => rst,
      outs_valid => source11_outs_valid,
      outs_ready => source11_outs_ready
    );

  constant50 : entity work.handshake_constant_3(arch) generic map(5)
    port map(
      ctrl_valid => source11_outs_valid,
      ctrl_ready => source11_outs_ready,
      clk => clk,
      rst => rst,
      outs => constant50_outs,
      outs_valid => constant50_outs_valid,
      outs_ready => constant50_outs_ready
    );

  extsi59 : entity work.extsi(arch) generic map(5, 6)
    port map(
      ins => constant50_outs,
      ins_valid => constant50_outs_valid,
      ins_ready => constant50_outs_ready,
      clk => clk,
      rst => rst,
      outs => extsi59_outs,
      outs_valid => extsi59_outs_valid,
      outs_ready => extsi59_outs_ready
    );

  source12 : entity work.source(arch)
    port map(
      clk => clk,
      rst => rst,
      outs_valid => source12_outs_valid,
      outs_ready => source12_outs_ready
    );

  constant51 : entity work.handshake_constant_1(arch) generic map(2)
    port map(
      ctrl_valid => source12_outs_valid,
      ctrl_ready => source12_outs_ready,
      clk => clk,
      rst => rst,
      outs => constant51_outs,
      outs_valid => constant51_outs_valid,
      outs_ready => constant51_outs_ready
    );

  fork61 : entity work.handshake_fork(arch) generic map(2, 2)
    port map(
      ins => constant51_outs,
      ins_valid => constant51_outs_valid,
      ins_ready => constant51_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork61_outs_0,
      outs(1) => fork61_outs_1,
      outs_valid(0) => fork61_outs_0_valid,
      outs_valid(1) => fork61_outs_1_valid,
      outs_ready(0) => fork61_outs_0_ready,
      outs_ready(1) => fork61_outs_1_ready
    );

  extsi60 : entity work.extsi(arch) generic map(2, 6)
    port map(
      ins => buffer138_outs,
      ins_valid => buffer138_outs_valid,
      ins_ready => buffer138_outs_ready,
      clk => clk,
      rst => rst,
      outs => extsi60_outs,
      outs_valid => extsi60_outs_valid,
      outs_ready => extsi60_outs_ready
    );

  buffer138 : entity work.tfifo(arch) generic map(1, 2)
    port map(
      ins => fork61_outs_0,
      ins_valid => fork61_outs_0_valid,
      ins_ready => fork61_outs_0_ready,
      clk => clk,
      rst => rst,
      outs => buffer138_outs,
      outs_valid => buffer138_outs_valid,
      outs_ready => buffer138_outs_ready
    );

  extsi23 : entity work.extsi(arch) generic map(2, 32)
    port map(
      ins => buffer139_outs,
      ins_valid => buffer139_outs_valid,
      ins_ready => buffer139_outs_ready,
      clk => clk,
      rst => rst,
      outs => extsi23_outs,
      outs_valid => extsi23_outs_valid,
      outs_ready => extsi23_outs_ready
    );

  buffer139 : entity work.tfifo(arch) generic map(1, 2)
    port map(
      ins => fork61_outs_1,
      ins_valid => fork61_outs_1_valid,
      ins_ready => fork61_outs_1_ready,
      clk => clk,
      rst => rst,
      outs => buffer139_outs,
      outs_valid => buffer139_outs_valid,
      outs_ready => buffer139_outs_ready
    );

  fork62 : entity work.handshake_fork(arch) generic map(4, 32)
    port map(
      ins => extsi23_outs,
      ins_valid => extsi23_outs_valid,
      ins_ready => extsi23_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork62_outs_0,
      outs(1) => fork62_outs_1,
      outs(2) => fork62_outs_2,
      outs(3) => fork62_outs_3,
      outs_valid(0) => fork62_outs_0_valid,
      outs_valid(1) => fork62_outs_1_valid,
      outs_valid(2) => fork62_outs_2_valid,
      outs_valid(3) => fork62_outs_3_valid,
      outs_ready(0) => fork62_outs_0_ready,
      outs_ready(1) => fork62_outs_1_ready,
      outs_ready(2) => fork62_outs_2_ready,
      outs_ready(3) => fork62_outs_3_ready
    );

  source13 : entity work.source(arch)
    port map(
      clk => clk,
      rst => rst,
      outs_valid => source13_outs_valid,
      outs_ready => source13_outs_ready
    );

  constant52 : entity work.handshake_constant_2(arch) generic map(3)
    port map(
      ctrl_valid => source13_outs_valid,
      ctrl_ready => source13_outs_ready,
      clk => clk,
      rst => rst,
      outs => constant52_outs,
      outs_valid => constant52_outs_valid,
      outs_ready => constant52_outs_ready
    );

  extsi24 : entity work.extsi(arch) generic map(3, 32)
    port map(
      ins => constant52_outs,
      ins_valid => constant52_outs_valid,
      ins_ready => constant52_outs_ready,
      clk => clk,
      rst => rst,
      outs => extsi24_outs,
      outs_valid => extsi24_outs_valid,
      outs_ready => extsi24_outs_ready
    );

  fork63 : entity work.handshake_fork(arch) generic map(4, 32)
    port map(
      ins => extsi24_outs,
      ins_valid => extsi24_outs_valid,
      ins_ready => extsi24_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork63_outs_0,
      outs(1) => fork63_outs_1,
      outs(2) => fork63_outs_2,
      outs(3) => fork63_outs_3,
      outs_valid(0) => fork63_outs_0_valid,
      outs_valid(1) => fork63_outs_1_valid,
      outs_valid(2) => fork63_outs_2_valid,
      outs_valid(3) => fork63_outs_3_valid,
      outs_ready(0) => fork63_outs_0_ready,
      outs_ready(1) => fork63_outs_1_ready,
      outs_ready(2) => fork63_outs_2_ready,
      outs_ready(3) => fork63_outs_3_ready
    );

  shli14 : entity work.shli(arch) generic map(32)
    port map(
      lhs => buffer141_outs,
      lhs_valid => buffer141_outs_valid,
      lhs_ready => buffer141_outs_ready,
      rhs => fork62_outs_0,
      rhs_valid => fork62_outs_0_valid,
      rhs_ready => fork62_outs_0_ready,
      clk => clk,
      rst => rst,
      result => shli14_result,
      result_valid => shli14_result_valid,
      result_ready => shli14_result_ready
    );

  buffer141 : entity work.tfifo(arch) generic map(1, 32)
    port map(
      ins => fork56_outs_0,
      ins_valid => fork56_outs_0_valid,
      ins_ready => fork56_outs_0_ready,
      clk => clk,
      rst => rst,
      outs => buffer141_outs,
      outs_valid => buffer141_outs_valid,
      outs_ready => buffer141_outs_ready
    );

  shli15 : entity work.shli(arch) generic map(32)
    port map(
      lhs => buffer143_outs,
      lhs_valid => buffer143_outs_valid,
      lhs_ready => buffer143_outs_ready,
      rhs => fork63_outs_0,
      rhs_valid => fork63_outs_0_valid,
      rhs_ready => fork63_outs_0_ready,
      clk => clk,
      rst => rst,
      result => shli15_result,
      result_valid => shli15_result_valid,
      result_ready => shli15_result_ready
    );

  buffer143 : entity work.tfifo(arch) generic map(1, 32)
    port map(
      ins => fork56_outs_1,
      ins_valid => fork56_outs_1_valid,
      ins_ready => fork56_outs_1_ready,
      clk => clk,
      rst => rst,
      outs => buffer143_outs,
      outs_valid => buffer143_outs_valid,
      outs_ready => buffer143_outs_ready
    );

  buffer197 : entity work.oehb(arch) generic map(32)
    port map(
      ins => shli14_result,
      ins_valid => shli14_result_valid,
      ins_ready => shli14_result_ready,
      clk => clk,
      rst => rst,
      outs => buffer197_outs,
      outs_valid => buffer197_outs_valid,
      outs_ready => buffer197_outs_ready
    );

  buffer198 : entity work.oehb(arch) generic map(32)
    port map(
      ins => shli15_result,
      ins_valid => shli15_result_valid,
      ins_ready => shli15_result_ready,
      clk => clk,
      rst => rst,
      outs => buffer198_outs,
      outs_valid => buffer198_outs_valid,
      outs_ready => buffer198_outs_ready
    );

  addi26 : entity work.addi(arch) generic map(32)
    port map(
      lhs => buffer197_outs,
      lhs_valid => buffer197_outs_valid,
      lhs_ready => buffer197_outs_ready,
      rhs => buffer198_outs,
      rhs_valid => buffer198_outs_valid,
      rhs_ready => buffer198_outs_ready,
      clk => clk,
      rst => rst,
      result => addi26_result,
      result_valid => addi26_result_valid,
      result_ready => addi26_result_ready
    );

  buffer199 : entity work.oehb(arch) generic map(32)
    port map(
      ins => addi26_result,
      ins_valid => addi26_result_valid,
      ins_ready => addi26_result_ready,
      clk => clk,
      rst => rst,
      outs => buffer199_outs,
      outs_valid => buffer199_outs_valid,
      outs_ready => buffer199_outs_ready
    );

  addi9 : entity work.addi(arch) generic map(32)
    port map(
      lhs => buffer144_outs,
      lhs_valid => buffer144_outs_valid,
      lhs_ready => buffer144_outs_ready,
      rhs => buffer199_outs,
      rhs_valid => buffer199_outs_valid,
      rhs_ready => buffer199_outs_ready,
      clk => clk,
      rst => rst,
      result => addi9_result,
      result_valid => addi9_result_valid,
      result_ready => addi9_result_ready
    );

  buffer144 : entity work.tfifo(arch) generic map(1, 32)
    port map(
      ins => fork54_outs_0,
      ins_valid => fork54_outs_0_valid,
      ins_ready => fork54_outs_0_ready,
      clk => clk,
      rst => rst,
      outs => buffer144_outs,
      outs_valid => buffer144_outs_valid,
      outs_ready => buffer144_outs_ready
    );

  gate2 : entity work.gate(arch) generic map(3, 32)
    port map(
      ins(0) => addi9_result,
      ins_valid(0) => addi9_result_valid,
      ins_valid(1) => fork51_outs_0_valid,
      ins_valid(2) => fork50_outs_0_valid,
      ins_ready(0) => addi9_result_ready,
      ins_ready(1) => fork51_outs_0_ready,
      ins_ready(2) => fork50_outs_0_ready,
      clk => clk,
      rst => rst,
      outs => gate2_outs,
      outs_valid => gate2_outs_valid,
      outs_ready => gate2_outs_ready
    );

  trunci15 : entity work.trunci(arch) generic map(32, 7)
    port map(
      ins => gate2_outs,
      ins_valid => gate2_outs_valid,
      ins_ready => gate2_outs_ready,
      clk => clk,
      rst => rst,
      outs => trunci15_outs,
      outs_valid => trunci15_outs_valid,
      outs_ready => trunci15_outs_ready
    );

  load4 : entity work.load(arch) generic map(32, 7)
    port map(
      addrIn => trunci15_outs,
      addrIn_valid => trunci15_outs_valid,
      addrIn_ready => trunci15_outs_ready,
      dataFromMem => mem_controller7_ldData_1,
      dataFromMem_valid => mem_controller7_ldData_1_valid,
      dataFromMem_ready => mem_controller7_ldData_1_ready,
      clk => clk,
      rst => rst,
      addrOut => load4_addrOut,
      addrOut_valid => load4_addrOut_valid,
      addrOut_ready => load4_addrOut_ready,
      dataOut => load4_dataOut,
      dataOut_valid => load4_dataOut_valid,
      dataOut_ready => load4_dataOut_ready
    );

  shli16 : entity work.shli(arch) generic map(32)
    port map(
      lhs => buffer146_outs,
      lhs_valid => buffer146_outs_valid,
      lhs_ready => buffer146_outs_ready,
      rhs => fork62_outs_1,
      rhs_valid => fork62_outs_1_valid,
      rhs_ready => fork62_outs_1_ready,
      clk => clk,
      rst => rst,
      result => shli16_result,
      result_valid => shli16_result_valid,
      result_ready => shli16_result_ready
    );

  buffer146 : entity work.tfifo(arch) generic map(1, 32)
    port map(
      ins => fork54_outs_1,
      ins_valid => fork54_outs_1_valid,
      ins_ready => fork54_outs_1_ready,
      clk => clk,
      rst => rst,
      outs => buffer146_outs,
      outs_valid => buffer146_outs_valid,
      outs_ready => buffer146_outs_ready
    );

  buffer200 : entity work.oehb(arch) generic map(32)
    port map(
      ins => shli16_result,
      ins_valid => shli16_result_valid,
      ins_ready => shli16_result_ready,
      clk => clk,
      rst => rst,
      outs => buffer200_outs,
      outs_valid => buffer200_outs_valid,
      outs_ready => buffer200_outs_ready
    );

  trunci16 : entity work.trunci(arch) generic map(32, 7)
    port map(
      ins => buffer200_outs,
      ins_valid => buffer200_outs_valid,
      ins_ready => buffer200_outs_ready,
      clk => clk,
      rst => rst,
      outs => trunci16_outs,
      outs_valid => trunci16_outs_valid,
      outs_ready => trunci16_outs_ready
    );

  shli17 : entity work.shli(arch) generic map(32)
    port map(
      lhs => buffer148_outs,
      lhs_valid => buffer148_outs_valid,
      lhs_ready => buffer148_outs_ready,
      rhs => fork63_outs_1,
      rhs_valid => fork63_outs_1_valid,
      rhs_ready => fork63_outs_1_ready,
      clk => clk,
      rst => rst,
      result => shli17_result,
      result_valid => shli17_result_valid,
      result_ready => shli17_result_ready
    );

  buffer148 : entity work.tfifo(arch) generic map(1, 32)
    port map(
      ins => fork54_outs_2,
      ins_valid => fork54_outs_2_valid,
      ins_ready => fork54_outs_2_ready,
      clk => clk,
      rst => rst,
      outs => buffer148_outs,
      outs_valid => buffer148_outs_valid,
      outs_ready => buffer148_outs_ready
    );

  buffer201 : entity work.oehb(arch) generic map(32)
    port map(
      ins => shli17_result,
      ins_valid => shli17_result_valid,
      ins_ready => shli17_result_ready,
      clk => clk,
      rst => rst,
      outs => buffer201_outs,
      outs_valid => buffer201_outs_valid,
      outs_ready => buffer201_outs_ready
    );

  trunci17 : entity work.trunci(arch) generic map(32, 7)
    port map(
      ins => buffer201_outs,
      ins_valid => buffer201_outs_valid,
      ins_ready => buffer201_outs_ready,
      clk => clk,
      rst => rst,
      outs => trunci17_outs,
      outs_valid => trunci17_outs_valid,
      outs_ready => trunci17_outs_ready
    );

  addi27 : entity work.addi(arch) generic map(7)
    port map(
      lhs => trunci16_outs,
      lhs_valid => trunci16_outs_valid,
      lhs_ready => trunci16_outs_ready,
      rhs => trunci17_outs,
      rhs_valid => trunci17_outs_valid,
      rhs_ready => trunci17_outs_ready,
      clk => clk,
      rst => rst,
      result => addi27_result,
      result_valid => addi27_result_valid,
      result_ready => addi27_result_ready
    );

  buffer202 : entity work.oehb(arch) generic map(7)
    port map(
      ins => addi27_result,
      ins_valid => addi27_result_valid,
      ins_ready => addi27_result_ready,
      clk => clk,
      rst => rst,
      outs => buffer202_outs,
      outs_valid => buffer202_outs_valid,
      outs_ready => buffer202_outs_ready
    );

  addi10 : entity work.addi(arch) generic map(7)
    port map(
      lhs => extsi57_outs,
      lhs_valid => extsi57_outs_valid,
      lhs_ready => extsi57_outs_ready,
      rhs => buffer202_outs,
      rhs_valid => buffer202_outs_valid,
      rhs_ready => buffer202_outs_ready,
      clk => clk,
      rst => rst,
      result => addi10_result,
      result_valid => addi10_result_valid,
      result_ready => addi10_result_ready
    );

  load5 : entity work.load(arch) generic map(32, 7)
    port map(
      addrIn => addi10_result,
      addrIn_valid => addi10_result_valid,
      addrIn_ready => addi10_result_ready,
      dataFromMem => mem_controller4_ldData_0,
      dataFromMem_valid => mem_controller4_ldData_0_valid,
      dataFromMem_ready => mem_controller4_ldData_0_ready,
      clk => clk,
      rst => rst,
      addrOut => load5_addrOut,
      addrOut_valid => load5_addrOut_valid,
      addrOut_ready => load5_addrOut_ready,
      dataOut => load5_dataOut,
      dataOut_valid => load5_dataOut_valid,
      dataOut_ready => load5_dataOut_ready
    );

  muli3 : entity work.muli(arch) generic map(32)
    port map(
      lhs => load4_dataOut,
      lhs_valid => load4_dataOut_valid,
      lhs_ready => load4_dataOut_ready,
      rhs => load5_dataOut,
      rhs_valid => load5_dataOut_valid,
      rhs_ready => load5_dataOut_ready,
      clk => clk,
      rst => rst,
      result => muli3_result,
      result_valid => muli3_result_valid,
      result_ready => muli3_result_ready
    );

  shli18 : entity work.shli(arch) generic map(32)
    port map(
      lhs => buffer150_outs,
      lhs_valid => buffer150_outs_valid,
      lhs_ready => buffer150_outs_ready,
      rhs => buffer149_outs,
      rhs_valid => buffer149_outs_valid,
      rhs_ready => buffer149_outs_ready,
      clk => clk,
      rst => rst,
      result => shli18_result,
      result_valid => shli18_result_valid,
      result_ready => shli18_result_ready
    );

  buffer149 : entity work.tfifo(arch) generic map(2, 32)
    port map(
      ins => fork62_outs_2,
      ins_valid => fork62_outs_2_valid,
      ins_ready => fork62_outs_2_ready,
      clk => clk,
      rst => rst,
      outs => buffer149_outs,
      outs_valid => buffer149_outs_valid,
      outs_ready => buffer149_outs_ready
    );

  buffer150 : entity work.tfifo(arch) generic map(2, 32)
    port map(
      ins => fork56_outs_2,
      ins_valid => fork56_outs_2_valid,
      ins_ready => fork56_outs_2_ready,
      clk => clk,
      rst => rst,
      outs => buffer150_outs,
      outs_valid => buffer150_outs_valid,
      outs_ready => buffer150_outs_ready
    );

  shli19 : entity work.shli(arch) generic map(32)
    port map(
      lhs => buffer152_outs,
      lhs_valid => buffer152_outs_valid,
      lhs_ready => buffer152_outs_ready,
      rhs => buffer151_outs,
      rhs_valid => buffer151_outs_valid,
      rhs_ready => buffer151_outs_ready,
      clk => clk,
      rst => rst,
      result => shli19_result,
      result_valid => shli19_result_valid,
      result_ready => shli19_result_ready
    );

  buffer151 : entity work.tfifo(arch) generic map(2, 32)
    port map(
      ins => fork63_outs_2,
      ins_valid => fork63_outs_2_valid,
      ins_ready => fork63_outs_2_ready,
      clk => clk,
      rst => rst,
      outs => buffer151_outs,
      outs_valid => buffer151_outs_valid,
      outs_ready => buffer151_outs_ready
    );

  buffer152 : entity work.tfifo(arch) generic map(2, 32)
    port map(
      ins => fork56_outs_3,
      ins_valid => fork56_outs_3_valid,
      ins_ready => fork56_outs_3_ready,
      clk => clk,
      rst => rst,
      outs => buffer152_outs,
      outs_valid => buffer152_outs_valid,
      outs_ready => buffer152_outs_ready
    );

  buffer203 : entity work.oehb(arch) generic map(32)
    port map(
      ins => shli18_result,
      ins_valid => shli18_result_valid,
      ins_ready => shli18_result_ready,
      clk => clk,
      rst => rst,
      outs => buffer203_outs,
      outs_valid => buffer203_outs_valid,
      outs_ready => buffer203_outs_ready
    );

  buffer204 : entity work.oehb(arch) generic map(32)
    port map(
      ins => shli19_result,
      ins_valid => shli19_result_valid,
      ins_ready => shli19_result_ready,
      clk => clk,
      rst => rst,
      outs => buffer204_outs,
      outs_valid => buffer204_outs_valid,
      outs_ready => buffer204_outs_ready
    );

  addi28 : entity work.addi(arch) generic map(32)
    port map(
      lhs => buffer203_outs,
      lhs_valid => buffer203_outs_valid,
      lhs_ready => buffer203_outs_ready,
      rhs => buffer204_outs,
      rhs_valid => buffer204_outs_valid,
      rhs_ready => buffer204_outs_ready,
      clk => clk,
      rst => rst,
      result => addi28_result,
      result_valid => addi28_result_valid,
      result_ready => addi28_result_ready
    );

  buffer205 : entity work.oehb(arch) generic map(32)
    port map(
      ins => addi28_result,
      ins_valid => addi28_result_valid,
      ins_ready => addi28_result_ready,
      clk => clk,
      rst => rst,
      outs => buffer205_outs,
      outs_valid => buffer205_outs_valid,
      outs_ready => buffer205_outs_ready
    );

  addi11 : entity work.addi(arch) generic map(32)
    port map(
      lhs => buffer153_outs,
      lhs_valid => buffer153_outs_valid,
      lhs_ready => buffer153_outs_ready,
      rhs => buffer205_outs,
      rhs_valid => buffer205_outs_valid,
      rhs_ready => buffer205_outs_ready,
      clk => clk,
      rst => rst,
      result => addi11_result,
      result_valid => addi11_result_valid,
      result_ready => addi11_result_ready
    );

  buffer153 : entity work.tfifo(arch) generic map(2, 32)
    port map(
      ins => fork58_outs_0,
      ins_valid => fork58_outs_0_valid,
      ins_ready => fork58_outs_0_ready,
      clk => clk,
      rst => rst,
      outs => buffer153_outs,
      outs_valid => buffer153_outs_valid,
      outs_ready => buffer153_outs_ready
    );

  buffer187 : entity work.tehb_dataless(arch)
    port map(
      ins_valid => mux52_outs_valid,
      ins_ready => mux52_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer187_outs_valid,
      outs_ready => buffer187_outs_ready
    );

  gate3 : entity work.gate(arch) generic map(3, 32)
    port map(
      ins(0) => addi11_result,
      ins_valid(0) => addi11_result_valid,
      ins_valid(1) => buffer187_outs_valid,
      ins_valid(2) => fork49_outs_1_valid,
      ins_ready(0) => addi11_result_ready,
      ins_ready(1) => buffer187_outs_ready,
      ins_ready(2) => fork49_outs_1_ready,
      clk => clk,
      rst => rst,
      outs => gate3_outs,
      outs_valid => gate3_outs_valid,
      outs_ready => gate3_outs_ready
    );

  trunci18 : entity work.trunci(arch) generic map(32, 7)
    port map(
      ins => gate3_outs,
      ins_valid => gate3_outs_valid,
      ins_ready => gate3_outs_ready,
      clk => clk,
      rst => rst,
      outs => trunci18_outs,
      outs_valid => trunci18_outs_valid,
      outs_ready => trunci18_outs_ready
    );

  load6 : entity work.load(arch) generic map(32, 7)
    port map(
      addrIn => trunci18_outs,
      addrIn_valid => trunci18_outs_valid,
      addrIn_ready => trunci18_outs_ready,
      dataFromMem => mem_controller3_ldData_1,
      dataFromMem_valid => mem_controller3_ldData_1_valid,
      dataFromMem_ready => mem_controller3_ldData_1_ready,
      clk => clk,
      rst => rst,
      addrOut => load6_addrOut,
      addrOut_valid => load6_addrOut_valid,
      addrOut_ready => load6_addrOut_ready,
      dataOut => load6_dataOut,
      dataOut_valid => load6_dataOut_valid,
      dataOut_ready => load6_dataOut_ready
    );

  addi1 : entity work.addi(arch) generic map(32)
    port map(
      lhs => load6_dataOut,
      lhs_valid => load6_dataOut_valid,
      lhs_ready => load6_dataOut_ready,
      rhs => muli3_result,
      rhs_valid => muli3_result_valid,
      rhs_ready => muli3_result_ready,
      clk => clk,
      rst => rst,
      result => addi1_result,
      result_valid => addi1_result_valid,
      result_ready => addi1_result_ready
    );

  shli20 : entity work.shli(arch) generic map(32)
    port map(
      lhs => buffer155_outs,
      lhs_valid => buffer155_outs_valid,
      lhs_ready => buffer155_outs_ready,
      rhs => buffer154_outs,
      rhs_valid => buffer154_outs_valid,
      rhs_ready => buffer154_outs_ready,
      clk => clk,
      rst => rst,
      result => shli20_result,
      result_valid => shli20_result_valid,
      result_ready => shli20_result_ready
    );

  buffer154 : entity work.tfifo(arch) generic map(3, 32)
    port map(
      ins => fork62_outs_3,
      ins_valid => fork62_outs_3_valid,
      ins_ready => fork62_outs_3_ready,
      clk => clk,
      rst => rst,
      outs => buffer154_outs,
      outs_valid => buffer154_outs_valid,
      outs_ready => buffer154_outs_ready
    );

  buffer155 : entity work.tfifo(arch) generic map(3, 32)
    port map(
      ins => fork56_outs_4,
      ins_valid => fork56_outs_4_valid,
      ins_ready => fork56_outs_4_ready,
      clk => clk,
      rst => rst,
      outs => buffer155_outs,
      outs_valid => buffer155_outs_valid,
      outs_ready => buffer155_outs_ready
    );

  shli21 : entity work.shli(arch) generic map(32)
    port map(
      lhs => buffer157_outs,
      lhs_valid => buffer157_outs_valid,
      lhs_ready => buffer157_outs_ready,
      rhs => buffer156_outs,
      rhs_valid => buffer156_outs_valid,
      rhs_ready => buffer156_outs_ready,
      clk => clk,
      rst => rst,
      result => shli21_result,
      result_valid => shli21_result_valid,
      result_ready => shli21_result_ready
    );

  buffer156 : entity work.tfifo(arch) generic map(3, 32)
    port map(
      ins => fork63_outs_3,
      ins_valid => fork63_outs_3_valid,
      ins_ready => fork63_outs_3_ready,
      clk => clk,
      rst => rst,
      outs => buffer156_outs,
      outs_valid => buffer156_outs_valid,
      outs_ready => buffer156_outs_ready
    );

  buffer157 : entity work.tfifo(arch) generic map(3, 32)
    port map(
      ins => fork56_outs_5,
      ins_valid => fork56_outs_5_valid,
      ins_ready => fork56_outs_5_ready,
      clk => clk,
      rst => rst,
      outs => buffer157_outs,
      outs_valid => buffer157_outs_valid,
      outs_ready => buffer157_outs_ready
    );

  buffer206 : entity work.oehb(arch) generic map(32)
    port map(
      ins => shli20_result,
      ins_valid => shli20_result_valid,
      ins_ready => shli20_result_ready,
      clk => clk,
      rst => rst,
      outs => buffer206_outs,
      outs_valid => buffer206_outs_valid,
      outs_ready => buffer206_outs_ready
    );

  buffer207 : entity work.oehb(arch) generic map(32)
    port map(
      ins => shli21_result,
      ins_valid => shli21_result_valid,
      ins_ready => shli21_result_ready,
      clk => clk,
      rst => rst,
      outs => buffer207_outs,
      outs_valid => buffer207_outs_valid,
      outs_ready => buffer207_outs_ready
    );

  addi29 : entity work.addi(arch) generic map(32)
    port map(
      lhs => buffer206_outs,
      lhs_valid => buffer206_outs_valid,
      lhs_ready => buffer206_outs_ready,
      rhs => buffer207_outs,
      rhs_valid => buffer207_outs_valid,
      rhs_ready => buffer207_outs_ready,
      clk => clk,
      rst => rst,
      result => addi29_result,
      result_valid => addi29_result_valid,
      result_ready => addi29_result_ready
    );

  buffer208 : entity work.oehb(arch) generic map(32)
    port map(
      ins => addi29_result,
      ins_valid => addi29_result_valid,
      ins_ready => addi29_result_ready,
      clk => clk,
      rst => rst,
      outs => buffer208_outs,
      outs_valid => buffer208_outs_valid,
      outs_ready => buffer208_outs_ready
    );

  addi12 : entity work.addi(arch) generic map(32)
    port map(
      lhs => buffer158_outs,
      lhs_valid => buffer158_outs_valid,
      lhs_ready => buffer158_outs_ready,
      rhs => buffer208_outs,
      rhs_valid => buffer208_outs_valid,
      rhs_ready => buffer208_outs_ready,
      clk => clk,
      rst => rst,
      result => addi12_result,
      result_valid => addi12_result_valid,
      result_ready => addi12_result_ready
    );

  buffer158 : entity work.tfifo(arch) generic map(2, 32)
    port map(
      ins => fork58_outs_1,
      ins_valid => fork58_outs_1_valid,
      ins_ready => fork58_outs_1_ready,
      clk => clk,
      rst => rst,
      outs => buffer158_outs,
      outs_valid => buffer158_outs_valid,
      outs_ready => buffer158_outs_ready
    );

  buffer4 : entity work.tfifo_dataless(arch) generic map(1)
    port map(
      ins_valid => store3_doneOut_valid,
      ins_ready => store3_doneOut_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer4_outs_valid,
      outs_ready => buffer4_outs_ready
    );

  gate4 : entity work.gate(arch) generic map(3, 32)
    port map(
      ins(0) => addi12_result,
      ins_valid(0) => addi12_result_valid,
      ins_valid(1) => fork52_outs_0_valid,
      ins_valid(2) => fork49_outs_0_valid,
      ins_ready(0) => addi12_result_ready,
      ins_ready(1) => fork52_outs_0_ready,
      ins_ready(2) => fork49_outs_0_ready,
      clk => clk,
      rst => rst,
      outs => gate4_outs,
      outs_valid => gate4_outs_valid,
      outs_ready => gate4_outs_ready
    );

  trunci19 : entity work.trunci(arch) generic map(32, 7)
    port map(
      ins => gate4_outs,
      ins_valid => gate4_outs_valid,
      ins_ready => gate4_outs_ready,
      clk => clk,
      rst => rst,
      outs => trunci19_outs,
      outs_valid => trunci19_outs_valid,
      outs_ready => trunci19_outs_ready
    );

  store3 : entity work.store(arch) generic map(32, 7)
    port map(
      addrIn => trunci19_outs,
      addrIn_valid => trunci19_outs_valid,
      addrIn_ready => trunci19_outs_ready,
      dataIn => addi1_result,
      dataIn_valid => addi1_result_valid,
      dataIn_ready => addi1_result_ready,
      doneFromMem_valid => mem_controller3_stDone_1_valid,
      doneFromMem_ready => mem_controller3_stDone_1_ready,
      clk => clk,
      rst => rst,
      addrOut => store3_addrOut,
      addrOut_valid => store3_addrOut_valid,
      addrOut_ready => store3_addrOut_ready,
      dataToMem => store3_dataToMem,
      dataToMem_valid => store3_dataToMem_valid,
      dataToMem_ready => store3_dataToMem_ready,
      doneOut_valid => store3_doneOut_valid,
      doneOut_ready => store3_doneOut_ready
    );

  addi16 : entity work.addi(arch) generic map(6)
    port map(
      lhs => extsi54_outs,
      lhs_valid => extsi54_outs_valid,
      lhs_ready => extsi54_outs_ready,
      rhs => extsi60_outs,
      rhs_valid => extsi60_outs_valid,
      rhs_ready => extsi60_outs_ready,
      clk => clk,
      rst => rst,
      result => addi16_result,
      result_valid => addi16_result_valid,
      result_ready => addi16_result_ready
    );

  fork64 : entity work.handshake_fork(arch) generic map(2, 6)
    port map(
      ins => addi16_result,
      ins_valid => addi16_result_valid,
      ins_ready => addi16_result_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork64_outs_0,
      outs(1) => fork64_outs_1,
      outs_valid(0) => fork64_outs_0_valid,
      outs_valid(1) => fork64_outs_1_valid,
      outs_ready(0) => fork64_outs_0_ready,
      outs_ready(1) => fork64_outs_1_ready
    );

  trunci20 : entity work.trunci(arch) generic map(6, 5)
    port map(
      ins => buffer159_outs,
      ins_valid => buffer159_outs_valid,
      ins_ready => buffer159_outs_ready,
      clk => clk,
      rst => rst,
      outs => trunci20_outs,
      outs_valid => trunci20_outs_valid,
      outs_ready => trunci20_outs_ready
    );

  buffer159 : entity work.tfifo(arch) generic map(1, 6)
    port map(
      ins => fork64_outs_0,
      ins_valid => fork64_outs_0_valid,
      ins_ready => fork64_outs_0_ready,
      clk => clk,
      rst => rst,
      outs => buffer159_outs,
      outs_valid => buffer159_outs_valid,
      outs_ready => buffer159_outs_ready
    );

  cmpi3 : entity work.handshake_cmpi_0(arch) generic map(6)
    port map(
      lhs => buffer160_outs,
      lhs_valid => buffer160_outs_valid,
      lhs_ready => buffer160_outs_ready,
      rhs => extsi59_outs,
      rhs_valid => extsi59_outs_valid,
      rhs_ready => extsi59_outs_ready,
      clk => clk,
      rst => rst,
      result => cmpi3_result,
      result_valid => cmpi3_result_valid,
      result_ready => cmpi3_result_ready
    );

  buffer210 : entity work.oehb(arch) generic map(6)
    port map(
      ins => fork64_outs_1,
      ins_valid => fork64_outs_1_valid,
      ins_ready => fork64_outs_1_ready,
      clk => clk,
      rst => rst,
      outs => buffer210_outs,
      outs_valid => buffer210_outs_valid,
      outs_ready => buffer210_outs_ready
    );

  buffer160 : entity work.tfifo(arch) generic map(1, 6)
    port map(
      ins => buffer210_outs,
      ins_valid => buffer210_outs_valid,
      ins_ready => buffer210_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer160_outs,
      outs_valid => buffer160_outs_valid,
      outs_ready => buffer160_outs_ready
    );

  buffer211 : entity work.oehb(arch) generic map(1)
    port map(
      ins => cmpi3_result,
      ins_valid => cmpi3_result_valid,
      ins_ready => cmpi3_result_ready,
      clk => clk,
      rst => rst,
      outs => buffer211_outs,
      outs_valid => buffer211_outs_valid,
      outs_ready => buffer211_outs_ready
    );

  fork65 : entity work.handshake_fork(arch) generic map(11, 1)
    port map(
      ins => buffer211_outs,
      ins_valid => buffer211_outs_valid,
      ins_ready => buffer211_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork65_outs_0,
      outs(1) => fork65_outs_1,
      outs(2) => fork65_outs_2,
      outs(3) => fork65_outs_3,
      outs(4) => fork65_outs_4,
      outs(5) => fork65_outs_5,
      outs(6) => fork65_outs_6,
      outs(7) => fork65_outs_7,
      outs(8) => fork65_outs_8,
      outs(9) => fork65_outs_9,
      outs(10) => fork65_outs_10,
      outs_valid(0) => fork65_outs_0_valid,
      outs_valid(1) => fork65_outs_1_valid,
      outs_valid(2) => fork65_outs_2_valid,
      outs_valid(3) => fork65_outs_3_valid,
      outs_valid(4) => fork65_outs_4_valid,
      outs_valid(5) => fork65_outs_5_valid,
      outs_valid(6) => fork65_outs_6_valid,
      outs_valid(7) => fork65_outs_7_valid,
      outs_valid(8) => fork65_outs_8_valid,
      outs_valid(9) => fork65_outs_9_valid,
      outs_valid(10) => fork65_outs_10_valid,
      outs_ready(0) => fork65_outs_0_ready,
      outs_ready(1) => fork65_outs_1_ready,
      outs_ready(2) => fork65_outs_2_ready,
      outs_ready(3) => fork65_outs_3_ready,
      outs_ready(4) => fork65_outs_4_ready,
      outs_ready(5) => fork65_outs_5_ready,
      outs_ready(6) => fork65_outs_6_ready,
      outs_ready(7) => fork65_outs_7_ready,
      outs_ready(8) => fork65_outs_8_ready,
      outs_ready(9) => fork65_outs_9_ready,
      outs_ready(10) => fork65_outs_10_ready
    );

  cond_br22 : entity work.cond_br(arch) generic map(5)
    port map(
      condition => fork65_outs_0,
      condition_valid => fork65_outs_0_valid,
      condition_ready => fork65_outs_0_ready,
      data => trunci20_outs,
      data_valid => trunci20_outs_valid,
      data_ready => trunci20_outs_ready,
      clk => clk,
      rst => rst,
      trueOut => cond_br22_trueOut,
      trueOut_valid => cond_br22_trueOut_valid,
      trueOut_ready => cond_br22_trueOut_ready,
      falseOut => cond_br22_falseOut,
      falseOut_valid => cond_br22_falseOut_valid,
      falseOut_ready => cond_br22_falseOut_ready
    );

  sink14 : entity work.sink(arch) generic map(5)
    port map(
      ins => cond_br22_falseOut,
      ins_valid => cond_br22_falseOut_valid,
      ins_ready => cond_br22_falseOut_ready,
      clk => clk,
      rst => rst
    );

  buffer190 : entity work.oehb(arch) generic map(32)
    port map(
      ins => mux18_outs,
      ins_valid => mux18_outs_valid,
      ins_ready => mux18_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer190_outs,
      outs_valid => buffer190_outs_valid,
      outs_ready => buffer190_outs_ready
    );

  buffer191 : entity work.tehb(arch) generic map(32)
    port map(
      ins => buffer190_outs,
      ins_valid => buffer190_outs_valid,
      ins_ready => buffer190_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer191_outs,
      outs_valid => buffer191_outs_valid,
      outs_ready => buffer191_outs_ready
    );

  cond_br23 : entity work.cond_br(arch) generic map(32)
    port map(
      condition => buffer162_outs,
      condition_valid => buffer162_outs_valid,
      condition_ready => buffer162_outs_ready,
      data => buffer191_outs,
      data_valid => buffer191_outs_valid,
      data_ready => buffer191_outs_ready,
      clk => clk,
      rst => rst,
      trueOut => cond_br23_trueOut,
      trueOut_valid => cond_br23_trueOut_valid,
      trueOut_ready => cond_br23_trueOut_ready,
      falseOut => cond_br23_falseOut,
      falseOut_valid => cond_br23_falseOut_valid,
      falseOut_ready => cond_br23_falseOut_ready
    );

  buffer162 : entity work.tfifo(arch) generic map(1, 1)
    port map(
      ins => fork65_outs_9,
      ins_valid => fork65_outs_9_valid,
      ins_ready => fork65_outs_9_ready,
      clk => clk,
      rst => rst,
      outs => buffer162_outs,
      outs_valid => buffer162_outs_valid,
      outs_ready => buffer162_outs_ready
    );

  cond_br24 : entity work.cond_br(arch) generic map(5)
    port map(
      condition => fork65_outs_1,
      condition_valid => fork65_outs_1_valid,
      condition_ready => fork65_outs_1_ready,
      data => buffer164_outs,
      data_valid => buffer164_outs_valid,
      data_ready => buffer164_outs_ready,
      clk => clk,
      rst => rst,
      trueOut => cond_br24_trueOut,
      trueOut_valid => cond_br24_trueOut_valid,
      trueOut_ready => cond_br24_trueOut_ready,
      falseOut => cond_br24_falseOut,
      falseOut_valid => cond_br24_falseOut_valid,
      falseOut_ready => cond_br24_falseOut_ready
    );

  buffer164 : entity work.tfifo(arch) generic map(1, 5)
    port map(
      ins => fork55_outs_0,
      ins_valid => fork55_outs_0_valid,
      ins_ready => fork55_outs_0_ready,
      clk => clk,
      rst => rst,
      outs => buffer164_outs,
      outs_valid => buffer164_outs_valid,
      outs_ready => buffer164_outs_ready
    );

  cond_br25 : entity work.cond_br(arch) generic map(5)
    port map(
      condition => fork65_outs_2,
      condition_valid => fork65_outs_2_valid,
      condition_ready => fork65_outs_2_ready,
      data => buffer166_outs,
      data_valid => buffer166_outs_valid,
      data_ready => buffer166_outs_ready,
      clk => clk,
      rst => rst,
      trueOut => cond_br25_trueOut,
      trueOut_valid => cond_br25_trueOut_valid,
      trueOut_ready => cond_br25_trueOut_ready,
      falseOut => cond_br25_falseOut,
      falseOut_valid => cond_br25_falseOut_valid,
      falseOut_ready => cond_br25_falseOut_ready
    );

  buffer166 : entity work.tfifo(arch) generic map(1, 5)
    port map(
      ins => fork57_outs_1,
      ins_valid => fork57_outs_1_valid,
      ins_ready => fork57_outs_1_ready,
      clk => clk,
      rst => rst,
      outs => buffer166_outs,
      outs_valid => buffer166_outs_valid,
      outs_ready => buffer166_outs_ready
    );

  cond_br26 : entity work.cond_br_dataless(arch)
    port map(
      condition => buffer167_outs,
      condition_valid => buffer167_outs_valid,
      condition_ready => buffer167_outs_ready,
      data_valid => fork60_outs_1_valid,
      data_ready => fork60_outs_1_ready,
      clk => clk,
      rst => rst,
      trueOut_valid => cond_br26_trueOut_valid,
      trueOut_ready => cond_br26_trueOut_ready,
      falseOut_valid => cond_br26_falseOut_valid,
      falseOut_ready => cond_br26_falseOut_ready
    );

  buffer167 : entity work.tfifo(arch) generic map(1, 1)
    port map(
      ins => fork65_outs_10,
      ins_valid => fork65_outs_10_valid,
      ins_ready => fork65_outs_10_ready,
      clk => clk,
      rst => rst,
      outs => buffer167_outs,
      outs_valid => buffer167_outs_valid,
      outs_ready => buffer167_outs_ready
    );

  cond_br94 : entity work.cond_br_dataless(arch)
    port map(
      condition => fork67_outs_4,
      condition_valid => fork67_outs_4_valid,
      condition_ready => fork67_outs_4_ready,
      data_valid => fork38_outs_0_valid,
      data_ready => fork38_outs_0_ready,
      clk => clk,
      rst => rst,
      trueOut_valid => cond_br94_trueOut_valid,
      trueOut_ready => cond_br94_trueOut_ready,
      falseOut_valid => cond_br94_falseOut_valid,
      falseOut_ready => cond_br94_falseOut_ready
    );

  sink15 : entity work.sink_dataless(arch)
    port map(
      ins_valid => cond_br94_falseOut_valid,
      ins_ready => cond_br94_falseOut_ready,
      clk => clk,
      rst => rst
    );

  cond_br95 : entity work.cond_br_dataless(arch)
    port map(
      condition => buffer169_outs,
      condition_valid => buffer169_outs_valid,
      condition_ready => buffer169_outs_ready,
      data_valid => fork37_outs_0_valid,
      data_ready => fork37_outs_0_ready,
      clk => clk,
      rst => rst,
      trueOut_valid => cond_br95_trueOut_valid,
      trueOut_ready => cond_br95_trueOut_ready,
      falseOut_valid => cond_br95_falseOut_valid,
      falseOut_ready => cond_br95_falseOut_ready
    );

  buffer169 : entity work.tfifo(arch) generic map(1, 1)
    port map(
      ins => fork67_outs_3,
      ins_valid => fork67_outs_3_valid,
      ins_ready => fork67_outs_3_ready,
      clk => clk,
      rst => rst,
      outs => buffer169_outs,
      outs_valid => buffer169_outs_valid,
      outs_ready => buffer169_outs_ready
    );

  sink16 : entity work.sink_dataless(arch)
    port map(
      ins_valid => cond_br95_falseOut_valid,
      ins_ready => cond_br95_falseOut_ready,
      clk => clk,
      rst => rst
    );

  cond_br96 : entity work.cond_br_dataless(arch)
    port map(
      condition => buffer170_outs,
      condition_valid => buffer170_outs_valid,
      condition_ready => buffer170_outs_ready,
      data_valid => cond_br93_falseOut_valid,
      data_ready => cond_br93_falseOut_ready,
      clk => clk,
      rst => rst,
      trueOut_valid => cond_br96_trueOut_valid,
      trueOut_ready => cond_br96_trueOut_ready,
      falseOut_valid => cond_br96_falseOut_valid,
      falseOut_ready => cond_br96_falseOut_ready
    );

  buffer170 : entity work.tfifo(arch) generic map(1, 1)
    port map(
      ins => fork67_outs_2,
      ins_valid => fork67_outs_2_valid,
      ins_ready => fork67_outs_2_ready,
      clk => clk,
      rst => rst,
      outs => buffer170_outs,
      outs_valid => buffer170_outs_valid,
      outs_ready => buffer170_outs_ready
    );

  extsi61 : entity work.extsi(arch) generic map(5, 6)
    port map(
      ins => cond_br25_falseOut,
      ins_valid => cond_br25_falseOut_valid,
      ins_ready => cond_br25_falseOut_ready,
      clk => clk,
      rst => rst,
      outs => extsi61_outs,
      outs_valid => extsi61_outs_valid,
      outs_ready => extsi61_outs_ready
    );

  source14 : entity work.source(arch)
    port map(
      clk => clk,
      rst => rst,
      outs_valid => source14_outs_valid,
      outs_ready => source14_outs_ready
    );

  constant53 : entity work.handshake_constant_3(arch) generic map(5)
    port map(
      ctrl_valid => source14_outs_valid,
      ctrl_ready => source14_outs_ready,
      clk => clk,
      rst => rst,
      outs => constant53_outs,
      outs_valid => constant53_outs_valid,
      outs_ready => constant53_outs_ready
    );

  extsi62 : entity work.extsi(arch) generic map(5, 6)
    port map(
      ins => constant53_outs,
      ins_valid => constant53_outs_valid,
      ins_ready => constant53_outs_ready,
      clk => clk,
      rst => rst,
      outs => extsi62_outs,
      outs_valid => extsi62_outs_valid,
      outs_ready => extsi62_outs_ready
    );

  source15 : entity work.source(arch)
    port map(
      clk => clk,
      rst => rst,
      outs_valid => source15_outs_valid,
      outs_ready => source15_outs_ready
    );

  constant54 : entity work.handshake_constant_1(arch) generic map(2)
    port map(
      ctrl_valid => source15_outs_valid,
      ctrl_ready => source15_outs_ready,
      clk => clk,
      rst => rst,
      outs => constant54_outs,
      outs_valid => constant54_outs_valid,
      outs_ready => constant54_outs_ready
    );

  extsi63 : entity work.extsi(arch) generic map(2, 6)
    port map(
      ins => constant54_outs,
      ins_valid => constant54_outs_valid,
      ins_ready => constant54_outs_ready,
      clk => clk,
      rst => rst,
      outs => extsi63_outs,
      outs_valid => extsi63_outs_valid,
      outs_ready => extsi63_outs_ready
    );

  addi17 : entity work.addi(arch) generic map(6)
    port map(
      lhs => extsi61_outs,
      lhs_valid => extsi61_outs_valid,
      lhs_ready => extsi61_outs_ready,
      rhs => extsi63_outs,
      rhs_valid => extsi63_outs_valid,
      rhs_ready => extsi63_outs_ready,
      clk => clk,
      rst => rst,
      result => addi17_result,
      result_valid => addi17_result_valid,
      result_ready => addi17_result_ready
    );

  buffer213 : entity work.oehb(arch) generic map(6)
    port map(
      ins => addi17_result,
      ins_valid => addi17_result_valid,
      ins_ready => addi17_result_ready,
      clk => clk,
      rst => rst,
      outs => buffer213_outs,
      outs_valid => buffer213_outs_valid,
      outs_ready => buffer213_outs_ready
    );

  fork66 : entity work.handshake_fork(arch) generic map(2, 6)
    port map(
      ins => buffer213_outs,
      ins_valid => buffer213_outs_valid,
      ins_ready => buffer213_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork66_outs_0,
      outs(1) => fork66_outs_1,
      outs_valid(0) => fork66_outs_0_valid,
      outs_valid(1) => fork66_outs_1_valid,
      outs_ready(0) => fork66_outs_0_ready,
      outs_ready(1) => fork66_outs_1_ready
    );

  trunci21 : entity work.trunci(arch) generic map(6, 5)
    port map(
      ins => fork66_outs_0,
      ins_valid => fork66_outs_0_valid,
      ins_ready => fork66_outs_0_ready,
      clk => clk,
      rst => rst,
      outs => trunci21_outs,
      outs_valid => trunci21_outs_valid,
      outs_ready => trunci21_outs_ready
    );

  cmpi4 : entity work.handshake_cmpi_0(arch) generic map(6)
    port map(
      lhs => fork66_outs_1,
      lhs_valid => fork66_outs_1_valid,
      lhs_ready => fork66_outs_1_ready,
      rhs => extsi62_outs,
      rhs_valid => extsi62_outs_valid,
      rhs_ready => extsi62_outs_ready,
      clk => clk,
      rst => rst,
      result => cmpi4_result,
      result_valid => cmpi4_result_valid,
      result_ready => cmpi4_result_ready
    );

  buffer214 : entity work.oehb(arch) generic map(1)
    port map(
      ins => cmpi4_result,
      ins_valid => cmpi4_result_valid,
      ins_ready => cmpi4_result_ready,
      clk => clk,
      rst => rst,
      outs => buffer214_outs,
      outs_valid => buffer214_outs_valid,
      outs_ready => buffer214_outs_ready
    );

  fork67 : entity work.handshake_fork(arch) generic map(8, 1)
    port map(
      ins => buffer214_outs,
      ins_valid => buffer214_outs_valid,
      ins_ready => buffer214_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork67_outs_0,
      outs(1) => fork67_outs_1,
      outs(2) => fork67_outs_2,
      outs(3) => fork67_outs_3,
      outs(4) => fork67_outs_4,
      outs(5) => fork67_outs_5,
      outs(6) => fork67_outs_6,
      outs(7) => fork67_outs_7,
      outs_valid(0) => fork67_outs_0_valid,
      outs_valid(1) => fork67_outs_1_valid,
      outs_valid(2) => fork67_outs_2_valid,
      outs_valid(3) => fork67_outs_3_valid,
      outs_valid(4) => fork67_outs_4_valid,
      outs_valid(5) => fork67_outs_5_valid,
      outs_valid(6) => fork67_outs_6_valid,
      outs_valid(7) => fork67_outs_7_valid,
      outs_ready(0) => fork67_outs_0_ready,
      outs_ready(1) => fork67_outs_1_ready,
      outs_ready(2) => fork67_outs_2_ready,
      outs_ready(3) => fork67_outs_3_ready,
      outs_ready(4) => fork67_outs_4_ready,
      outs_ready(5) => fork67_outs_5_ready,
      outs_ready(6) => fork67_outs_6_ready,
      outs_ready(7) => fork67_outs_7_ready
    );

  cond_br27 : entity work.cond_br(arch) generic map(5)
    port map(
      condition => fork67_outs_0,
      condition_valid => fork67_outs_0_valid,
      condition_ready => fork67_outs_0_ready,
      data => trunci21_outs,
      data_valid => trunci21_outs_valid,
      data_ready => trunci21_outs_ready,
      clk => clk,
      rst => rst,
      trueOut => cond_br27_trueOut,
      trueOut_valid => cond_br27_trueOut_valid,
      trueOut_ready => cond_br27_trueOut_ready,
      falseOut => cond_br27_falseOut,
      falseOut_valid => cond_br27_falseOut_valid,
      falseOut_ready => cond_br27_falseOut_ready
    );

  sink18 : entity work.sink(arch) generic map(5)
    port map(
      ins => cond_br27_falseOut,
      ins_valid => cond_br27_falseOut_valid,
      ins_ready => cond_br27_falseOut_ready,
      clk => clk,
      rst => rst
    );

  buffer212 : entity work.oehb(arch) generic map(32)
    port map(
      ins => cond_br23_falseOut,
      ins_valid => cond_br23_falseOut_valid,
      ins_ready => cond_br23_falseOut_ready,
      clk => clk,
      rst => rst,
      outs => buffer212_outs,
      outs_valid => buffer212_outs_valid,
      outs_ready => buffer212_outs_ready
    );

  cond_br28 : entity work.cond_br(arch) generic map(32)
    port map(
      condition => buffer174_outs,
      condition_valid => buffer174_outs_valid,
      condition_ready => buffer174_outs_ready,
      data => buffer212_outs,
      data_valid => buffer212_outs_valid,
      data_ready => buffer212_outs_ready,
      clk => clk,
      rst => rst,
      trueOut => cond_br28_trueOut,
      trueOut_valid => cond_br28_trueOut_valid,
      trueOut_ready => cond_br28_trueOut_ready,
      falseOut => cond_br28_falseOut,
      falseOut_valid => cond_br28_falseOut_valid,
      falseOut_ready => cond_br28_falseOut_ready
    );

  buffer174 : entity work.tfifo(arch) generic map(1, 1)
    port map(
      ins => fork67_outs_6,
      ins_valid => fork67_outs_6_valid,
      ins_ready => fork67_outs_6_ready,
      clk => clk,
      rst => rst,
      outs => buffer174_outs,
      outs_valid => buffer174_outs_valid,
      outs_ready => buffer174_outs_ready
    );

  cond_br29 : entity work.cond_br(arch) generic map(5)
    port map(
      condition => fork67_outs_1,
      condition_valid => fork67_outs_1_valid,
      condition_ready => fork67_outs_1_ready,
      data => cond_br24_falseOut,
      data_valid => cond_br24_falseOut_valid,
      data_ready => cond_br24_falseOut_ready,
      clk => clk,
      rst => rst,
      trueOut => cond_br29_trueOut,
      trueOut_valid => cond_br29_trueOut_valid,
      trueOut_ready => cond_br29_trueOut_ready,
      falseOut => cond_br29_falseOut,
      falseOut_valid => cond_br29_falseOut_valid,
      falseOut_ready => cond_br29_falseOut_ready
    );

  cond_br30 : entity work.cond_br_dataless(arch)
    port map(
      condition => buffer176_outs,
      condition_valid => buffer176_outs_valid,
      condition_ready => buffer176_outs_ready,
      data_valid => cond_br26_falseOut_valid,
      data_ready => cond_br26_falseOut_ready,
      clk => clk,
      rst => rst,
      trueOut_valid => cond_br30_trueOut_valid,
      trueOut_ready => cond_br30_trueOut_ready,
      falseOut_valid => cond_br30_falseOut_valid,
      falseOut_ready => cond_br30_falseOut_ready
    );

  buffer176 : entity work.tfifo(arch) generic map(1, 1)
    port map(
      ins => fork67_outs_7,
      ins_valid => fork67_outs_7_valid,
      ins_ready => fork67_outs_7_ready,
      clk => clk,
      rst => rst,
      outs => buffer176_outs,
      outs_valid => buffer176_outs_valid,
      outs_ready => buffer176_outs_ready
    );

  cond_br97 : entity work.cond_br_dataless(arch)
    port map(
      condition => buffer177_outs,
      condition_valid => buffer177_outs_valid,
      condition_ready => buffer177_outs_ready,
      data_valid => cond_br96_falseOut_valid,
      data_ready => cond_br96_falseOut_ready,
      clk => clk,
      rst => rst,
      trueOut_valid => cond_br97_trueOut_valid,
      trueOut_ready => cond_br97_trueOut_ready,
      falseOut_valid => cond_br97_falseOut_valid,
      falseOut_ready => cond_br97_falseOut_ready
    );

  buffer177 : entity work.tfifo(arch) generic map(1, 1)
    port map(
      ins => fork69_outs_3,
      ins_valid => fork69_outs_3_valid,
      ins_ready => fork69_outs_3_ready,
      clk => clk,
      rst => rst,
      outs => buffer177_outs,
      outs_valid => buffer177_outs_valid,
      outs_ready => buffer177_outs_ready
    );

  sink19 : entity work.sink_dataless(arch)
    port map(
      ins_valid => cond_br97_falseOut_valid,
      ins_ready => cond_br97_falseOut_ready,
      clk => clk,
      rst => rst
    );

  cond_br98 : entity work.cond_br_dataless(arch)
    port map(
      condition => fork69_outs_2,
      condition_valid => fork69_outs_2_valid,
      condition_ready => fork69_outs_2_ready,
      data_valid => fork33_outs_0_valid,
      data_ready => fork33_outs_0_ready,
      clk => clk,
      rst => rst,
      trueOut_valid => cond_br98_trueOut_valid,
      trueOut_ready => cond_br98_trueOut_ready,
      falseOut_valid => cond_br98_falseOut_valid,
      falseOut_ready => cond_br98_falseOut_ready
    );

  sink20 : entity work.sink_dataless(arch)
    port map(
      ins_valid => cond_br98_falseOut_valid,
      ins_ready => cond_br98_falseOut_ready,
      clk => clk,
      rst => rst
    );

  cond_br99 : entity work.cond_br_dataless(arch)
    port map(
      condition => fork69_outs_1,
      condition_valid => fork69_outs_1_valid,
      condition_ready => fork69_outs_1_ready,
      data_valid => fork32_outs_0_valid,
      data_ready => fork32_outs_0_ready,
      clk => clk,
      rst => rst,
      trueOut_valid => cond_br99_trueOut_valid,
      trueOut_ready => cond_br99_trueOut_ready,
      falseOut_valid => cond_br99_falseOut_valid,
      falseOut_ready => cond_br99_falseOut_ready
    );

  sink21 : entity work.sink_dataless(arch)
    port map(
      ins_valid => cond_br99_falseOut_valid,
      ins_ready => cond_br99_falseOut_ready,
      clk => clk,
      rst => rst
    );

  extsi64 : entity work.extsi(arch) generic map(5, 6)
    port map(
      ins => cond_br29_falseOut,
      ins_valid => cond_br29_falseOut_valid,
      ins_ready => cond_br29_falseOut_ready,
      clk => clk,
      rst => rst,
      outs => extsi64_outs,
      outs_valid => extsi64_outs_valid,
      outs_ready => extsi64_outs_ready
    );

  source16 : entity work.source(arch)
    port map(
      clk => clk,
      rst => rst,
      outs_valid => source16_outs_valid,
      outs_ready => source16_outs_ready
    );

  constant55 : entity work.handshake_constant_3(arch) generic map(5)
    port map(
      ctrl_valid => source16_outs_valid,
      ctrl_ready => source16_outs_ready,
      clk => clk,
      rst => rst,
      outs => constant55_outs,
      outs_valid => constant55_outs_valid,
      outs_ready => constant55_outs_ready
    );

  extsi65 : entity work.extsi(arch) generic map(5, 6)
    port map(
      ins => constant55_outs,
      ins_valid => constant55_outs_valid,
      ins_ready => constant55_outs_ready,
      clk => clk,
      rst => rst,
      outs => extsi65_outs,
      outs_valid => extsi65_outs_valid,
      outs_ready => extsi65_outs_ready
    );

  source17 : entity work.source(arch)
    port map(
      clk => clk,
      rst => rst,
      outs_valid => source17_outs_valid,
      outs_ready => source17_outs_ready
    );

  constant56 : entity work.handshake_constant_1(arch) generic map(2)
    port map(
      ctrl_valid => source17_outs_valid,
      ctrl_ready => source17_outs_ready,
      clk => clk,
      rst => rst,
      outs => constant56_outs,
      outs_valid => constant56_outs_valid,
      outs_ready => constant56_outs_ready
    );

  extsi66 : entity work.extsi(arch) generic map(2, 6)
    port map(
      ins => constant56_outs,
      ins_valid => constant56_outs_valid,
      ins_ready => constant56_outs_ready,
      clk => clk,
      rst => rst,
      outs => extsi66_outs,
      outs_valid => extsi66_outs_valid,
      outs_ready => extsi66_outs_ready
    );

  buffer216 : entity work.oehb(arch) generic map(6)
    port map(
      ins => extsi64_outs,
      ins_valid => extsi64_outs_valid,
      ins_ready => extsi64_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer216_outs,
      outs_valid => buffer216_outs_valid,
      outs_ready => buffer216_outs_ready
    );

  addi18 : entity work.addi(arch) generic map(6)
    port map(
      lhs => buffer216_outs,
      lhs_valid => buffer216_outs_valid,
      lhs_ready => buffer216_outs_ready,
      rhs => extsi66_outs,
      rhs_valid => extsi66_outs_valid,
      rhs_ready => extsi66_outs_ready,
      clk => clk,
      rst => rst,
      result => addi18_result,
      result_valid => addi18_result_valid,
      result_ready => addi18_result_ready
    );

  buffer217 : entity work.oehb(arch) generic map(6)
    port map(
      ins => addi18_result,
      ins_valid => addi18_result_valid,
      ins_ready => addi18_result_ready,
      clk => clk,
      rst => rst,
      outs => buffer217_outs,
      outs_valid => buffer217_outs_valid,
      outs_ready => buffer217_outs_ready
    );

  fork68 : entity work.handshake_fork(arch) generic map(2, 6)
    port map(
      ins => buffer217_outs,
      ins_valid => buffer217_outs_valid,
      ins_ready => buffer217_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork68_outs_0,
      outs(1) => fork68_outs_1,
      outs_valid(0) => fork68_outs_0_valid,
      outs_valid(1) => fork68_outs_1_valid,
      outs_ready(0) => fork68_outs_0_ready,
      outs_ready(1) => fork68_outs_1_ready
    );

  trunci22 : entity work.trunci(arch) generic map(6, 5)
    port map(
      ins => fork68_outs_0,
      ins_valid => fork68_outs_0_valid,
      ins_ready => fork68_outs_0_ready,
      clk => clk,
      rst => rst,
      outs => trunci22_outs,
      outs_valid => trunci22_outs_valid,
      outs_ready => trunci22_outs_ready
    );

  cmpi5 : entity work.handshake_cmpi_0(arch) generic map(6)
    port map(
      lhs => fork68_outs_1,
      lhs_valid => fork68_outs_1_valid,
      lhs_ready => fork68_outs_1_ready,
      rhs => extsi65_outs,
      rhs_valid => extsi65_outs_valid,
      rhs_ready => extsi65_outs_ready,
      clk => clk,
      rst => rst,
      result => cmpi5_result,
      result_valid => cmpi5_result_valid,
      result_ready => cmpi5_result_ready
    );

  buffer218 : entity work.oehb(arch) generic map(1)
    port map(
      ins => cmpi5_result,
      ins_valid => cmpi5_result_valid,
      ins_ready => cmpi5_result_ready,
      clk => clk,
      rst => rst,
      outs => buffer218_outs,
      outs_valid => buffer218_outs_valid,
      outs_ready => buffer218_outs_ready
    );

  fork69 : entity work.handshake_fork(arch) generic map(7, 1)
    port map(
      ins => buffer218_outs,
      ins_valid => buffer218_outs_valid,
      ins_ready => buffer218_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork69_outs_0,
      outs(1) => fork69_outs_1,
      outs(2) => fork69_outs_2,
      outs(3) => fork69_outs_3,
      outs(4) => fork69_outs_4,
      outs(5) => fork69_outs_5,
      outs(6) => fork69_outs_6,
      outs_valid(0) => fork69_outs_0_valid,
      outs_valid(1) => fork69_outs_1_valid,
      outs_valid(2) => fork69_outs_2_valid,
      outs_valid(3) => fork69_outs_3_valid,
      outs_valid(4) => fork69_outs_4_valid,
      outs_valid(5) => fork69_outs_5_valid,
      outs_valid(6) => fork69_outs_6_valid,
      outs_ready(0) => fork69_outs_0_ready,
      outs_ready(1) => fork69_outs_1_ready,
      outs_ready(2) => fork69_outs_2_ready,
      outs_ready(3) => fork69_outs_3_ready,
      outs_ready(4) => fork69_outs_4_ready,
      outs_ready(5) => fork69_outs_5_ready,
      outs_ready(6) => fork69_outs_6_ready
    );

  cond_br31 : entity work.cond_br(arch) generic map(5)
    port map(
      condition => fork69_outs_0,
      condition_valid => fork69_outs_0_valid,
      condition_ready => fork69_outs_0_ready,
      data => trunci22_outs,
      data_valid => trunci22_outs_valid,
      data_ready => trunci22_outs_ready,
      clk => clk,
      rst => rst,
      trueOut => cond_br31_trueOut,
      trueOut_valid => cond_br31_trueOut_valid,
      trueOut_ready => cond_br31_trueOut_ready,
      falseOut => cond_br31_falseOut,
      falseOut_valid => cond_br31_falseOut_valid,
      falseOut_ready => cond_br31_falseOut_ready
    );

  sink23 : entity work.sink(arch) generic map(5)
    port map(
      ins => cond_br31_falseOut,
      ins_valid => cond_br31_falseOut_valid,
      ins_ready => cond_br31_falseOut_ready,
      clk => clk,
      rst => rst
    );

  cond_br32 : entity work.cond_br(arch) generic map(32)
    port map(
      condition => fork69_outs_5,
      condition_valid => fork69_outs_5_valid,
      condition_ready => fork69_outs_5_ready,
      data => cond_br28_falseOut,
      data_valid => cond_br28_falseOut_valid,
      data_ready => cond_br28_falseOut_ready,
      clk => clk,
      rst => rst,
      trueOut => cond_br32_trueOut,
      trueOut_valid => cond_br32_trueOut_valid,
      trueOut_ready => cond_br32_trueOut_ready,
      falseOut => cond_br32_falseOut,
      falseOut_valid => cond_br32_falseOut_valid,
      falseOut_ready => cond_br32_falseOut_ready
    );

  sink24 : entity work.sink(arch) generic map(32)
    port map(
      ins => cond_br32_falseOut,
      ins_valid => cond_br32_falseOut_valid,
      ins_ready => cond_br32_falseOut_ready,
      clk => clk,
      rst => rst
    );

  cond_br33 : entity work.cond_br_dataless(arch)
    port map(
      condition => buffer184_outs,
      condition_valid => buffer184_outs_valid,
      condition_ready => buffer184_outs_ready,
      data_valid => cond_br30_falseOut_valid,
      data_ready => cond_br30_falseOut_ready,
      clk => clk,
      rst => rst,
      trueOut_valid => cond_br33_trueOut_valid,
      trueOut_ready => cond_br33_trueOut_ready,
      falseOut_valid => cond_br33_falseOut_valid,
      falseOut_ready => cond_br33_falseOut_ready
    );

  buffer184 : entity work.tfifo(arch) generic map(1, 1)
    port map(
      ins => fork69_outs_6,
      ins_valid => fork69_outs_6_valid,
      ins_ready => fork69_outs_6_ready,
      clk => clk,
      rst => rst,
      outs => buffer184_outs,
      outs_valid => buffer184_outs_valid,
      outs_ready => buffer184_outs_ready
    );

  fork70 : entity work.fork_dataless(arch) generic map(5)
    port map(
      ins_valid => cond_br33_falseOut_valid,
      ins_ready => cond_br33_falseOut_ready,
      clk => clk,
      rst => rst,
      outs_valid(0) => fork70_outs_0_valid,
      outs_valid(1) => fork70_outs_1_valid,
      outs_valid(2) => fork70_outs_2_valid,
      outs_valid(3) => fork70_outs_3_valid,
      outs_valid(4) => fork70_outs_4_valid,
      outs_ready(0) => fork70_outs_0_ready,
      outs_ready(1) => fork70_outs_1_ready,
      outs_ready(2) => fork70_outs_2_ready,
      outs_ready(3) => fork70_outs_3_ready,
      outs_ready(4) => fork70_outs_4_ready
    );

end architecture;
