library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity tfifo is
  generic (
    SIZE     : integer;
    BITWIDTH : integer
  );
  port (
    -- inputs
    clk, rst   : in std_logic;
    ins        : in std_logic_vector(BITWIDTH - 1 downto 0);
    ins_valid  : in std_logic;
    outs_ready : in std_logic;
    -- outputs
    outs       : out std_logic_vector(BITWIDTH - 1 downto 0);
    outs_valid : out std_logic
    outs_ready : out std_logic;
  );
end entity;

architecture arch of tfifo is
  signal mux_sel : std_logic;
  signal fifo_valid, fifo_ready : std_logic;
  signal fifo_pvalid, fifo_nready : std_logic;
  signal fifo_in, fifo_out : std_logic_vector(BITWIDTH - 1 downto 0);
begin

  process (mux_sel, fifo_out, ins) is
  begin
    if (mux_sel = '1') then
      outs <= fifo_out;
    else
      outs <= ins;
    end if;
  end process;

  outs_valid <= ins_valid or fifo_valid;
  outs_ready <= fifo_ready or outs_ready;
  fifo_pvalid <= ins_valid and (not outs_ready or fifo_valid);
  mux_sel <= fifo_valid;

  fifo_nready <= outs_ready;
  fifo_in <= ins;

  fifo : entity work.elastic_fifo_inner(arch) generic map (SIZE, BITWIDTH)
    port map(
      -- inputs
      clk        => clk,
      rst        => rst,
      ins        => fifo_in,
      ins_valid  => fifo_pvalid,
      outs_ready => fifo_nready,
      -- outputs
      outs       => fifo_out,
      outs_valid => fifo_valid,
      ins_ready  => fifo_ready,
    );

end arch;
