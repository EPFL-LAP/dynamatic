library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity bicg is
  port (
    q_loadData : in std_logic_vector(31 downto 0);
    q_start_valid : in std_logic;
    start_valid : in std_logic;
    clk : in std_logic;
    rst : in std_logic;
    out0_ready : in std_logic;
    q_end_ready : in std_logic;
    end_ready : in std_logic;
    q_start_ready : out std_logic;
    start_ready : out std_logic;
    out0 : out std_logic_vector(31 downto 0);
    out0_valid : out std_logic;
    q_end_valid : out std_logic;
    end_valid : out std_logic;
    q_loadEn : out std_logic;
    q_loadAddr : out std_logic_vector(4 downto 0);
    q_storeEn : out std_logic;
    q_storeAddr : out std_logic_vector(4 downto 0);
    q_storeData : out std_logic_vector(31 downto 0)
  );
end entity;

architecture behavioral of bicg is

  signal fork0_outs_0_valid : std_logic;
  signal fork0_outs_0_ready : std_logic;
  signal fork0_outs_1_valid : std_logic;
  signal fork0_outs_1_ready : std_logic;
  signal fork0_outs_2_valid : std_logic;
  signal fork0_outs_2_ready : std_logic;
  signal fork0_outs_3_valid : std_logic;
  signal fork0_outs_3_ready : std_logic;
  signal fork0_outs_4_valid : std_logic;
  signal fork0_outs_4_ready : std_logic;
  signal buffer20_outs_valid : std_logic;
  signal buffer20_outs_ready : std_logic;
  signal buffer21_outs_valid : std_logic;
  signal buffer21_outs_ready : std_logic;
  signal buffer22_outs_valid : std_logic;
  signal buffer22_outs_ready : std_logic;
  signal buffer23_outs_valid : std_logic;
  signal buffer23_outs_ready : std_logic;
  signal buffer24_outs_valid : std_logic;
  signal buffer24_outs_ready : std_logic;
  signal mem_controller1_memEnd_valid : std_logic;
  signal mem_controller1_memEnd_ready : std_logic;
  signal mem_controller1_loadEn : std_logic;
  signal mem_controller1_loadAddr : std_logic_vector(4 downto 0);
  signal mem_controller1_storeEn : std_logic;
  signal mem_controller1_storeAddr : std_logic_vector(4 downto 0);
  signal mem_controller1_storeData : std_logic_vector(31 downto 0);
  signal buffer15_outs_valid : std_logic;
  signal buffer15_outs_ready : std_logic;
  signal buffer16_outs_valid : std_logic;
  signal buffer16_outs_ready : std_logic;
  signal buffer17_outs_valid : std_logic;
  signal buffer17_outs_ready : std_logic;
  signal buffer18_outs_valid : std_logic;
  signal buffer18_outs_ready : std_logic;
  signal buffer19_outs_valid : std_logic;
  signal buffer19_outs_ready : std_logic;
  signal constant0_outs : std_logic_vector(0 downto 0);
  signal constant0_outs_valid : std_logic;
  signal constant0_outs_ready : std_logic;
  signal fork1_outs_0 : std_logic_vector(0 downto 0);
  signal fork1_outs_0_valid : std_logic;
  signal fork1_outs_0_ready : std_logic;
  signal fork1_outs_1 : std_logic_vector(0 downto 0);
  signal fork1_outs_1_valid : std_logic;
  signal fork1_outs_1_ready : std_logic;
  signal buffer30_outs : std_logic_vector(0 downto 0);
  signal buffer30_outs_valid : std_logic;
  signal buffer30_outs_ready : std_logic;
  signal buffer31_outs : std_logic_vector(0 downto 0);
  signal buffer31_outs_valid : std_logic;
  signal buffer31_outs_ready : std_logic;
  signal buffer32_outs : std_logic_vector(0 downto 0);
  signal buffer32_outs_valid : std_logic;
  signal buffer32_outs_ready : std_logic;
  signal buffer33_outs : std_logic_vector(0 downto 0);
  signal buffer33_outs_valid : std_logic;
  signal buffer33_outs_ready : std_logic;
  signal buffer34_outs : std_logic_vector(0 downto 0);
  signal buffer34_outs_valid : std_logic;
  signal buffer34_outs_ready : std_logic;
  signal extsi7_outs : std_logic_vector(5 downto 0);
  signal extsi7_outs_valid : std_logic;
  signal extsi7_outs_ready : std_logic;
  signal buffer25_outs : std_logic_vector(0 downto 0);
  signal buffer25_outs_valid : std_logic;
  signal buffer25_outs_ready : std_logic;
  signal buffer26_outs : std_logic_vector(0 downto 0);
  signal buffer26_outs_valid : std_logic;
  signal buffer26_outs_ready : std_logic;
  signal buffer27_outs : std_logic_vector(0 downto 0);
  signal buffer27_outs_valid : std_logic;
  signal buffer27_outs_ready : std_logic;
  signal buffer28_outs : std_logic_vector(0 downto 0);
  signal buffer28_outs_valid : std_logic;
  signal buffer28_outs_ready : std_logic;
  signal buffer29_outs : std_logic_vector(0 downto 0);
  signal buffer29_outs_valid : std_logic;
  signal buffer29_outs_ready : std_logic;
  signal buffer196_outs : std_logic_vector(0 downto 0);
  signal buffer196_outs_valid : std_logic;
  signal buffer196_outs_ready : std_logic;
  signal buffer197_outs : std_logic_vector(0 downto 0);
  signal buffer197_outs_valid : std_logic;
  signal buffer197_outs_ready : std_logic;
  signal buffer198_outs : std_logic_vector(0 downto 0);
  signal buffer198_outs_valid : std_logic;
  signal buffer198_outs_ready : std_logic;
  signal buffer199_outs : std_logic_vector(0 downto 0);
  signal buffer199_outs_valid : std_logic;
  signal buffer199_outs_ready : std_logic;
  signal buffer200_outs : std_logic_vector(0 downto 0);
  signal buffer200_outs_valid : std_logic;
  signal buffer200_outs_ready : std_logic;
  signal merge0_outs : std_logic_vector(0 downto 0);
  signal merge0_outs_valid : std_logic;
  signal merge0_outs_ready : std_logic;
  signal buffer35_outs : std_logic_vector(0 downto 0);
  signal buffer35_outs_valid : std_logic;
  signal buffer35_outs_ready : std_logic;
  signal fork2_outs_0 : std_logic_vector(0 downto 0);
  signal fork2_outs_0_valid : std_logic;
  signal fork2_outs_0_ready : std_logic;
  signal fork2_outs_1 : std_logic_vector(0 downto 0);
  signal fork2_outs_1_valid : std_logic;
  signal fork2_outs_1_ready : std_logic;
  signal buffer10_outs_valid : std_logic;
  signal buffer10_outs_ready : std_logic;
  signal buffer11_outs_valid : std_logic;
  signal buffer11_outs_ready : std_logic;
  signal buffer12_outs_valid : std_logic;
  signal buffer12_outs_ready : std_logic;
  signal buffer13_outs_valid : std_logic;
  signal buffer13_outs_ready : std_logic;
  signal buffer14_outs_valid : std_logic;
  signal buffer14_outs_ready : std_logic;
  signal buffer41_outs : std_logic_vector(0 downto 0);
  signal buffer41_outs_valid : std_logic;
  signal buffer41_outs_ready : std_logic;
  signal buffer42_outs : std_logic_vector(0 downto 0);
  signal buffer42_outs_valid : std_logic;
  signal buffer42_outs_ready : std_logic;
  signal buffer43_outs : std_logic_vector(0 downto 0);
  signal buffer43_outs_valid : std_logic;
  signal buffer43_outs_ready : std_logic;
  signal buffer44_outs : std_logic_vector(0 downto 0);
  signal buffer44_outs_valid : std_logic;
  signal buffer44_outs_ready : std_logic;
  signal buffer45_outs : std_logic_vector(0 downto 0);
  signal buffer45_outs_valid : std_logic;
  signal buffer45_outs_ready : std_logic;
  signal mux0_outs_valid : std_logic;
  signal mux0_outs_ready : std_logic;
  signal buffer46_outs_valid : std_logic;
  signal buffer46_outs_ready : std_logic;
  signal buffer47_outs_valid : std_logic;
  signal buffer47_outs_ready : std_logic;
  signal buffer48_outs_valid : std_logic;
  signal buffer48_outs_ready : std_logic;
  signal buffer49_outs_valid : std_logic;
  signal buffer49_outs_ready : std_logic;
  signal buffer50_outs_valid : std_logic;
  signal buffer50_outs_ready : std_logic;
  signal buffer51_outs_valid : std_logic;
  signal buffer51_outs_ready : std_logic;
  signal fork3_outs_0_valid : std_logic;
  signal fork3_outs_0_ready : std_logic;
  signal fork3_outs_1_valid : std_logic;
  signal fork3_outs_1_ready : std_logic;
  signal fork3_outs_2_valid : std_logic;
  signal fork3_outs_2_ready : std_logic;
  signal fork3_outs_3_valid : std_logic;
  signal fork3_outs_3_ready : std_logic;
  signal fork3_outs_4_valid : std_logic;
  signal fork3_outs_4_ready : std_logic;
  signal buffer36_outs : std_logic_vector(0 downto 0);
  signal buffer36_outs_valid : std_logic;
  signal buffer36_outs_ready : std_logic;
  signal buffer37_outs : std_logic_vector(0 downto 0);
  signal buffer37_outs_valid : std_logic;
  signal buffer37_outs_ready : std_logic;
  signal buffer38_outs : std_logic_vector(0 downto 0);
  signal buffer38_outs_valid : std_logic;
  signal buffer38_outs_ready : std_logic;
  signal buffer39_outs : std_logic_vector(0 downto 0);
  signal buffer39_outs_valid : std_logic;
  signal buffer39_outs_ready : std_logic;
  signal buffer40_outs : std_logic_vector(0 downto 0);
  signal buffer40_outs_valid : std_logic;
  signal buffer40_outs_ready : std_logic;
  signal mux5_outs : std_logic_vector(5 downto 0);
  signal mux5_outs_valid : std_logic;
  signal mux5_outs_ready : std_logic;
  signal buffer77_outs : std_logic_vector(5 downto 0);
  signal buffer77_outs_valid : std_logic;
  signal buffer77_outs_ready : std_logic;
  signal buffer78_outs : std_logic_vector(5 downto 0);
  signal buffer78_outs_valid : std_logic;
  signal buffer78_outs_ready : std_logic;
  signal buffer79_outs : std_logic_vector(5 downto 0);
  signal buffer79_outs_valid : std_logic;
  signal buffer79_outs_ready : std_logic;
  signal buffer80_outs : std_logic_vector(5 downto 0);
  signal buffer80_outs_valid : std_logic;
  signal buffer80_outs_ready : std_logic;
  signal buffer81_outs : std_logic_vector(5 downto 0);
  signal buffer81_outs_valid : std_logic;
  signal buffer81_outs_ready : std_logic;
  signal buffer82_outs : std_logic_vector(5 downto 0);
  signal buffer82_outs_valid : std_logic;
  signal buffer82_outs_ready : std_logic;
  signal fork4_outs_0 : std_logic_vector(5 downto 0);
  signal fork4_outs_0_valid : std_logic;
  signal fork4_outs_0_ready : std_logic;
  signal fork4_outs_1 : std_logic_vector(5 downto 0);
  signal fork4_outs_1_valid : std_logic;
  signal fork4_outs_1_ready : std_logic;
  signal fork4_outs_2 : std_logic_vector(5 downto 0);
  signal fork4_outs_2_valid : std_logic;
  signal fork4_outs_2_ready : std_logic;
  signal buffer93_outs : std_logic_vector(5 downto 0);
  signal buffer93_outs_valid : std_logic;
  signal buffer93_outs_ready : std_logic;
  signal buffer94_outs : std_logic_vector(5 downto 0);
  signal buffer94_outs_valid : std_logic;
  signal buffer94_outs_ready : std_logic;
  signal buffer95_outs : std_logic_vector(5 downto 0);
  signal buffer95_outs_valid : std_logic;
  signal buffer95_outs_ready : std_logic;
  signal buffer96_outs : std_logic_vector(5 downto 0);
  signal buffer96_outs_valid : std_logic;
  signal buffer96_outs_ready : std_logic;
  signal buffer97_outs : std_logic_vector(5 downto 0);
  signal buffer97_outs_valid : std_logic;
  signal buffer97_outs_ready : std_logic;
  signal extsi8_outs : std_logic_vector(6 downto 0);
  signal extsi8_outs_valid : std_logic;
  signal extsi8_outs_ready : std_logic;
  signal buffer88_outs : std_logic_vector(5 downto 0);
  signal buffer88_outs_valid : std_logic;
  signal buffer88_outs_ready : std_logic;
  signal buffer89_outs : std_logic_vector(5 downto 0);
  signal buffer89_outs_valid : std_logic;
  signal buffer89_outs_ready : std_logic;
  signal buffer90_outs : std_logic_vector(5 downto 0);
  signal buffer90_outs_valid : std_logic;
  signal buffer90_outs_ready : std_logic;
  signal buffer91_outs : std_logic_vector(5 downto 0);
  signal buffer91_outs_valid : std_logic;
  signal buffer91_outs_ready : std_logic;
  signal buffer92_outs : std_logic_vector(5 downto 0);
  signal buffer92_outs_valid : std_logic;
  signal buffer92_outs_ready : std_logic;
  signal extsi9_outs : std_logic_vector(31 downto 0);
  signal extsi9_outs_valid : std_logic;
  signal extsi9_outs_ready : std_logic;
  signal buffer83_outs : std_logic_vector(5 downto 0);
  signal buffer83_outs_valid : std_logic;
  signal buffer83_outs_ready : std_logic;
  signal buffer84_outs : std_logic_vector(5 downto 0);
  signal buffer84_outs_valid : std_logic;
  signal buffer84_outs_ready : std_logic;
  signal buffer85_outs : std_logic_vector(5 downto 0);
  signal buffer85_outs_valid : std_logic;
  signal buffer85_outs_ready : std_logic;
  signal buffer86_outs : std_logic_vector(5 downto 0);
  signal buffer86_outs_valid : std_logic;
  signal buffer86_outs_ready : std_logic;
  signal buffer87_outs : std_logic_vector(5 downto 0);
  signal buffer87_outs_valid : std_logic;
  signal buffer87_outs_ready : std_logic;
  signal trunci0_outs : std_logic_vector(4 downto 0);
  signal trunci0_outs_valid : std_logic;
  signal trunci0_outs_ready : std_logic;
  signal buffer72_outs_valid : std_logic;
  signal buffer72_outs_ready : std_logic;
  signal buffer73_outs_valid : std_logic;
  signal buffer73_outs_ready : std_logic;
  signal buffer74_outs_valid : std_logic;
  signal buffer74_outs_ready : std_logic;
  signal buffer75_outs_valid : std_logic;
  signal buffer75_outs_ready : std_logic;
  signal buffer76_outs_valid : std_logic;
  signal buffer76_outs_ready : std_logic;
  signal constant8_outs : std_logic_vector(0 downto 0);
  signal constant8_outs_valid : std_logic;
  signal constant8_outs_ready : std_logic;
  signal extsi10_outs : std_logic_vector(5 downto 0);
  signal extsi10_outs_valid : std_logic;
  signal extsi10_outs_ready : std_logic;
  signal buffer171_outs : std_logic_vector(0 downto 0);
  signal buffer171_outs_valid : std_logic;
  signal buffer171_outs_ready : std_logic;
  signal buffer172_outs : std_logic_vector(0 downto 0);
  signal buffer172_outs_valid : std_logic;
  signal buffer172_outs_ready : std_logic;
  signal buffer173_outs : std_logic_vector(0 downto 0);
  signal buffer173_outs_valid : std_logic;
  signal buffer173_outs_ready : std_logic;
  signal buffer174_outs : std_logic_vector(0 downto 0);
  signal buffer174_outs_valid : std_logic;
  signal buffer174_outs_ready : std_logic;
  signal buffer175_outs : std_logic_vector(0 downto 0);
  signal buffer175_outs_valid : std_logic;
  signal buffer175_outs_ready : std_logic;
  signal cond_br17_trueOut : std_logic_vector(31 downto 0);
  signal cond_br17_trueOut_valid : std_logic;
  signal cond_br17_trueOut_ready : std_logic;
  signal cond_br17_falseOut : std_logic_vector(31 downto 0);
  signal cond_br17_falseOut_valid : std_logic;
  signal cond_br17_falseOut_ready : std_logic;
  signal fork5_outs_0 : std_logic_vector(31 downto 0);
  signal fork5_outs_0_valid : std_logic;
  signal fork5_outs_0_ready : std_logic;
  signal fork5_outs_1 : std_logic_vector(31 downto 0);
  signal fork5_outs_1_valid : std_logic;
  signal fork5_outs_1_ready : std_logic;
  signal buffer176_outs : std_logic_vector(0 downto 0);
  signal buffer176_outs_valid : std_logic;
  signal buffer176_outs_ready : std_logic;
  signal buffer177_outs : std_logic_vector(0 downto 0);
  signal buffer177_outs_valid : std_logic;
  signal buffer177_outs_ready : std_logic;
  signal buffer178_outs : std_logic_vector(0 downto 0);
  signal buffer178_outs_valid : std_logic;
  signal buffer178_outs_ready : std_logic;
  signal buffer179_outs : std_logic_vector(0 downto 0);
  signal buffer179_outs_valid : std_logic;
  signal buffer179_outs_ready : std_logic;
  signal buffer180_outs : std_logic_vector(0 downto 0);
  signal buffer180_outs_valid : std_logic;
  signal buffer180_outs_ready : std_logic;
  signal cond_br18_trueOut : std_logic_vector(5 downto 0);
  signal cond_br18_trueOut_valid : std_logic;
  signal cond_br18_trueOut_ready : std_logic;
  signal cond_br18_falseOut : std_logic_vector(5 downto 0);
  signal cond_br18_falseOut_valid : std_logic;
  signal cond_br18_falseOut_ready : std_logic;
  signal buffer134_outs_valid : std_logic;
  signal buffer134_outs_ready : std_logic;
  signal buffer135_outs_valid : std_logic;
  signal buffer135_outs_ready : std_logic;
  signal buffer136_outs_valid : std_logic;
  signal buffer136_outs_ready : std_logic;
  signal buffer137_outs_valid : std_logic;
  signal buffer137_outs_ready : std_logic;
  signal buffer138_outs_valid : std_logic;
  signal buffer138_outs_ready : std_logic;
  signal buffer181_outs : std_logic_vector(0 downto 0);
  signal buffer181_outs_valid : std_logic;
  signal buffer181_outs_ready : std_logic;
  signal buffer182_outs : std_logic_vector(0 downto 0);
  signal buffer182_outs_valid : std_logic;
  signal buffer182_outs_ready : std_logic;
  signal buffer183_outs : std_logic_vector(0 downto 0);
  signal buffer183_outs_valid : std_logic;
  signal buffer183_outs_ready : std_logic;
  signal buffer184_outs : std_logic_vector(0 downto 0);
  signal buffer184_outs_valid : std_logic;
  signal buffer184_outs_ready : std_logic;
  signal buffer185_outs : std_logic_vector(0 downto 0);
  signal buffer185_outs_valid : std_logic;
  signal buffer185_outs_ready : std_logic;
  signal cond_br19_trueOut_valid : std_logic;
  signal cond_br19_trueOut_ready : std_logic;
  signal cond_br19_falseOut_valid : std_logic;
  signal cond_br19_falseOut_ready : std_logic;
  signal buffer67_outs_valid : std_logic;
  signal buffer67_outs_ready : std_logic;
  signal buffer68_outs_valid : std_logic;
  signal buffer68_outs_ready : std_logic;
  signal buffer69_outs_valid : std_logic;
  signal buffer69_outs_ready : std_logic;
  signal buffer70_outs_valid : std_logic;
  signal buffer70_outs_ready : std_logic;
  signal buffer71_outs_valid : std_logic;
  signal buffer71_outs_ready : std_logic;
  signal control_merge0_outs_valid : std_logic;
  signal control_merge0_outs_ready : std_logic;
  signal control_merge0_index : std_logic_vector(0 downto 0);
  signal control_merge0_index_valid : std_logic;
  signal control_merge0_index_ready : std_logic;
  signal fork6_outs_0 : std_logic_vector(0 downto 0);
  signal fork6_outs_0_valid : std_logic;
  signal fork6_outs_0_ready : std_logic;
  signal fork6_outs_1 : std_logic_vector(0 downto 0);
  signal fork6_outs_1_valid : std_logic;
  signal fork6_outs_1_ready : std_logic;
  signal buffer108_outs_valid : std_logic;
  signal buffer108_outs_ready : std_logic;
  signal buffer109_outs_valid : std_logic;
  signal buffer109_outs_ready : std_logic;
  signal buffer110_outs_valid : std_logic;
  signal buffer110_outs_ready : std_logic;
  signal buffer111_outs_valid : std_logic;
  signal buffer111_outs_ready : std_logic;
  signal buffer112_outs_valid : std_logic;
  signal buffer112_outs_ready : std_logic;
  signal buffer113_outs_valid : std_logic;
  signal buffer113_outs_ready : std_logic;
  signal fork7_outs_0_valid : std_logic;
  signal fork7_outs_0_ready : std_logic;
  signal fork7_outs_1_valid : std_logic;
  signal fork7_outs_1_ready : std_logic;
  signal fork7_outs_2_valid : std_logic;
  signal fork7_outs_2_ready : std_logic;
  signal buffer119_outs : std_logic_vector(0 downto 0);
  signal buffer119_outs_valid : std_logic;
  signal buffer119_outs_ready : std_logic;
  signal buffer120_outs : std_logic_vector(0 downto 0);
  signal buffer120_outs_valid : std_logic;
  signal buffer120_outs_ready : std_logic;
  signal buffer121_outs : std_logic_vector(0 downto 0);
  signal buffer121_outs_valid : std_logic;
  signal buffer121_outs_ready : std_logic;
  signal buffer122_outs : std_logic_vector(0 downto 0);
  signal buffer122_outs_valid : std_logic;
  signal buffer122_outs_ready : std_logic;
  signal buffer123_outs : std_logic_vector(0 downto 0);
  signal buffer123_outs_valid : std_logic;
  signal buffer123_outs_ready : std_logic;
  signal mux8_outs : std_logic_vector(31 downto 0);
  signal mux8_outs_valid : std_logic;
  signal mux8_outs_ready : std_logic;
  signal buffer114_outs : std_logic_vector(0 downto 0);
  signal buffer114_outs_valid : std_logic;
  signal buffer114_outs_ready : std_logic;
  signal buffer115_outs : std_logic_vector(0 downto 0);
  signal buffer115_outs_valid : std_logic;
  signal buffer115_outs_ready : std_logic;
  signal buffer116_outs : std_logic_vector(0 downto 0);
  signal buffer116_outs_valid : std_logic;
  signal buffer116_outs_ready : std_logic;
  signal buffer117_outs : std_logic_vector(0 downto 0);
  signal buffer117_outs_valid : std_logic;
  signal buffer117_outs_ready : std_logic;
  signal buffer118_outs : std_logic_vector(0 downto 0);
  signal buffer118_outs_valid : std_logic;
  signal buffer118_outs_ready : std_logic;
  signal mux9_outs : std_logic_vector(5 downto 0);
  signal mux9_outs_valid : std_logic;
  signal mux9_outs_ready : std_logic;
  signal buffer145_outs : std_logic_vector(5 downto 0);
  signal buffer145_outs_valid : std_logic;
  signal buffer145_outs_ready : std_logic;
  signal buffer146_outs : std_logic_vector(5 downto 0);
  signal buffer146_outs_valid : std_logic;
  signal buffer146_outs_ready : std_logic;
  signal buffer147_outs : std_logic_vector(5 downto 0);
  signal buffer147_outs_valid : std_logic;
  signal buffer147_outs_ready : std_logic;
  signal buffer148_outs : std_logic_vector(5 downto 0);
  signal buffer148_outs_valid : std_logic;
  signal buffer148_outs_ready : std_logic;
  signal buffer149_outs : std_logic_vector(5 downto 0);
  signal buffer149_outs_valid : std_logic;
  signal buffer149_outs_ready : std_logic;
  signal buffer150_outs : std_logic_vector(5 downto 0);
  signal buffer150_outs_valid : std_logic;
  signal buffer150_outs_ready : std_logic;
  signal fork8_outs_0 : std_logic_vector(5 downto 0);
  signal fork8_outs_0_valid : std_logic;
  signal fork8_outs_0_ready : std_logic;
  signal fork8_outs_1 : std_logic_vector(5 downto 0);
  signal fork8_outs_1_valid : std_logic;
  signal fork8_outs_1_ready : std_logic;
  signal buffer156_outs : std_logic_vector(5 downto 0);
  signal buffer156_outs_valid : std_logic;
  signal buffer156_outs_ready : std_logic;
  signal buffer157_outs : std_logic_vector(5 downto 0);
  signal buffer157_outs_valid : std_logic;
  signal buffer157_outs_ready : std_logic;
  signal buffer158_outs : std_logic_vector(5 downto 0);
  signal buffer158_outs_valid : std_logic;
  signal buffer158_outs_ready : std_logic;
  signal buffer159_outs : std_logic_vector(5 downto 0);
  signal buffer159_outs_valid : std_logic;
  signal buffer159_outs_ready : std_logic;
  signal buffer160_outs : std_logic_vector(5 downto 0);
  signal buffer160_outs_valid : std_logic;
  signal buffer160_outs_ready : std_logic;
  signal extsi11_outs : std_logic_vector(6 downto 0);
  signal extsi11_outs_valid : std_logic;
  signal extsi11_outs_ready : std_logic;
  signal buffer151_outs : std_logic_vector(5 downto 0);
  signal buffer151_outs_valid : std_logic;
  signal buffer151_outs_ready : std_logic;
  signal buffer152_outs : std_logic_vector(5 downto 0);
  signal buffer152_outs_valid : std_logic;
  signal buffer152_outs_ready : std_logic;
  signal buffer153_outs : std_logic_vector(5 downto 0);
  signal buffer153_outs_valid : std_logic;
  signal buffer153_outs_ready : std_logic;
  signal buffer154_outs : std_logic_vector(5 downto 0);
  signal buffer154_outs_valid : std_logic;
  signal buffer154_outs_ready : std_logic;
  signal buffer155_outs : std_logic_vector(5 downto 0);
  signal buffer155_outs_valid : std_logic;
  signal buffer155_outs_ready : std_logic;
  signal extsi12_outs : std_logic_vector(31 downto 0);
  signal extsi12_outs_valid : std_logic;
  signal extsi12_outs_ready : std_logic;
  signal buffer129_outs_valid : std_logic;
  signal buffer129_outs_ready : std_logic;
  signal buffer130_outs_valid : std_logic;
  signal buffer130_outs_ready : std_logic;
  signal buffer131_outs_valid : std_logic;
  signal buffer131_outs_ready : std_logic;
  signal buffer132_outs_valid : std_logic;
  signal buffer132_outs_ready : std_logic;
  signal buffer133_outs_valid : std_logic;
  signal buffer133_outs_ready : std_logic;
  signal constant9_outs : std_logic_vector(5 downto 0);
  signal constant9_outs_valid : std_logic;
  signal constant9_outs_ready : std_logic;
  signal extsi13_outs : std_logic_vector(6 downto 0);
  signal extsi13_outs_valid : std_logic;
  signal extsi13_outs_ready : std_logic;
  signal buffer124_outs_valid : std_logic;
  signal buffer124_outs_ready : std_logic;
  signal buffer125_outs_valid : std_logic;
  signal buffer125_outs_ready : std_logic;
  signal buffer126_outs_valid : std_logic;
  signal buffer126_outs_ready : std_logic;
  signal buffer127_outs_valid : std_logic;
  signal buffer127_outs_ready : std_logic;
  signal buffer128_outs_valid : std_logic;
  signal buffer128_outs_ready : std_logic;
  signal constant10_outs : std_logic_vector(1 downto 0);
  signal constant10_outs_valid : std_logic;
  signal constant10_outs_ready : std_logic;
  signal extsi14_outs : std_logic_vector(6 downto 0);
  signal extsi14_outs_valid : std_logic;
  signal extsi14_outs_ready : std_logic;
  signal buffer139_outs : std_logic_vector(31 downto 0);
  signal buffer139_outs_valid : std_logic;
  signal buffer139_outs_ready : std_logic;
  signal buffer140_outs : std_logic_vector(31 downto 0);
  signal buffer140_outs_valid : std_logic;
  signal buffer140_outs_ready : std_logic;
  signal buffer141_outs : std_logic_vector(31 downto 0);
  signal buffer141_outs_valid : std_logic;
  signal buffer141_outs_ready : std_logic;
  signal buffer142_outs : std_logic_vector(31 downto 0);
  signal buffer142_outs_valid : std_logic;
  signal buffer142_outs_ready : std_logic;
  signal buffer143_outs : std_logic_vector(31 downto 0);
  signal buffer143_outs_valid : std_logic;
  signal buffer143_outs_ready : std_logic;
  signal buffer144_outs : std_logic_vector(31 downto 0);
  signal buffer144_outs_valid : std_logic;
  signal buffer144_outs_ready : std_logic;
  signal muli0_result : std_logic_vector(31 downto 0);
  signal muli0_result_valid : std_logic;
  signal muli0_result_ready : std_logic;
  signal addi1_result : std_logic_vector(6 downto 0);
  signal addi1_result_valid : std_logic;
  signal addi1_result_ready : std_logic;
  signal fork9_outs_0 : std_logic_vector(6 downto 0);
  signal fork9_outs_0_valid : std_logic;
  signal fork9_outs_0_ready : std_logic;
  signal fork9_outs_1 : std_logic_vector(6 downto 0);
  signal fork9_outs_1_valid : std_logic;
  signal fork9_outs_1_ready : std_logic;
  signal buffer166_outs : std_logic_vector(6 downto 0);
  signal buffer166_outs_valid : std_logic;
  signal buffer166_outs_ready : std_logic;
  signal buffer167_outs : std_logic_vector(6 downto 0);
  signal buffer167_outs_valid : std_logic;
  signal buffer167_outs_ready : std_logic;
  signal buffer168_outs : std_logic_vector(6 downto 0);
  signal buffer168_outs_valid : std_logic;
  signal buffer168_outs_ready : std_logic;
  signal buffer169_outs : std_logic_vector(6 downto 0);
  signal buffer169_outs_valid : std_logic;
  signal buffer169_outs_ready : std_logic;
  signal buffer170_outs : std_logic_vector(6 downto 0);
  signal buffer170_outs_valid : std_logic;
  signal buffer170_outs_ready : std_logic;
  signal trunci1_outs : std_logic_vector(5 downto 0);
  signal trunci1_outs_valid : std_logic;
  signal trunci1_outs_ready : std_logic;
  signal buffer161_outs : std_logic_vector(6 downto 0);
  signal buffer161_outs_valid : std_logic;
  signal buffer161_outs_ready : std_logic;
  signal buffer162_outs : std_logic_vector(6 downto 0);
  signal buffer162_outs_valid : std_logic;
  signal buffer162_outs_ready : std_logic;
  signal buffer163_outs : std_logic_vector(6 downto 0);
  signal buffer163_outs_valid : std_logic;
  signal buffer163_outs_ready : std_logic;
  signal buffer164_outs : std_logic_vector(6 downto 0);
  signal buffer164_outs_valid : std_logic;
  signal buffer164_outs_ready : std_logic;
  signal buffer165_outs : std_logic_vector(6 downto 0);
  signal buffer165_outs_valid : std_logic;
  signal buffer165_outs_ready : std_logic;
  signal cmpi0_result : std_logic_vector(0 downto 0);
  signal cmpi0_result_valid : std_logic;
  signal cmpi0_result_ready : std_logic;
  signal fork10_outs_0 : std_logic_vector(0 downto 0);
  signal fork10_outs_0_valid : std_logic;
  signal fork10_outs_0_ready : std_logic;
  signal fork10_outs_1 : std_logic_vector(0 downto 0);
  signal fork10_outs_1_valid : std_logic;
  signal fork10_outs_1_ready : std_logic;
  signal fork10_outs_2 : std_logic_vector(0 downto 0);
  signal fork10_outs_2_valid : std_logic;
  signal fork10_outs_2_ready : std_logic;
  signal buffer103_outs : std_logic_vector(31 downto 0);
  signal buffer103_outs_valid : std_logic;
  signal buffer103_outs_ready : std_logic;
  signal buffer104_outs : std_logic_vector(31 downto 0);
  signal buffer104_outs_valid : std_logic;
  signal buffer104_outs_ready : std_logic;
  signal buffer105_outs : std_logic_vector(31 downto 0);
  signal buffer105_outs_valid : std_logic;
  signal buffer105_outs_ready : std_logic;
  signal buffer106_outs : std_logic_vector(31 downto 0);
  signal buffer106_outs_valid : std_logic;
  signal buffer106_outs_ready : std_logic;
  signal buffer107_outs : std_logic_vector(31 downto 0);
  signal buffer107_outs_valid : std_logic;
  signal buffer107_outs_ready : std_logic;
  signal buffer201_outs : std_logic_vector(0 downto 0);
  signal buffer201_outs_valid : std_logic;
  signal buffer201_outs_ready : std_logic;
  signal buffer202_outs : std_logic_vector(0 downto 0);
  signal buffer202_outs_valid : std_logic;
  signal buffer202_outs_ready : std_logic;
  signal buffer203_outs : std_logic_vector(0 downto 0);
  signal buffer203_outs_valid : std_logic;
  signal buffer203_outs_ready : std_logic;
  signal buffer204_outs : std_logic_vector(0 downto 0);
  signal buffer204_outs_valid : std_logic;
  signal buffer204_outs_ready : std_logic;
  signal buffer205_outs : std_logic_vector(0 downto 0);
  signal buffer205_outs_valid : std_logic;
  signal buffer205_outs_ready : std_logic;
  signal cond_br20_trueOut : std_logic_vector(31 downto 0);
  signal cond_br20_trueOut_valid : std_logic;
  signal cond_br20_trueOut_ready : std_logic;
  signal cond_br20_falseOut : std_logic_vector(31 downto 0);
  signal cond_br20_falseOut_valid : std_logic;
  signal cond_br20_falseOut_ready : std_logic;
  signal buffer206_outs : std_logic_vector(0 downto 0);
  signal buffer206_outs_valid : std_logic;
  signal buffer206_outs_ready : std_logic;
  signal buffer207_outs : std_logic_vector(0 downto 0);
  signal buffer207_outs_valid : std_logic;
  signal buffer207_outs_ready : std_logic;
  signal buffer208_outs : std_logic_vector(0 downto 0);
  signal buffer208_outs_valid : std_logic;
  signal buffer208_outs_ready : std_logic;
  signal buffer209_outs : std_logic_vector(0 downto 0);
  signal buffer209_outs_valid : std_logic;
  signal buffer209_outs_ready : std_logic;
  signal buffer210_outs : std_logic_vector(0 downto 0);
  signal buffer210_outs_valid : std_logic;
  signal buffer210_outs_ready : std_logic;
  signal cond_br21_trueOut : std_logic_vector(5 downto 0);
  signal cond_br21_trueOut_valid : std_logic;
  signal cond_br21_trueOut_ready : std_logic;
  signal cond_br21_falseOut : std_logic_vector(5 downto 0);
  signal cond_br21_falseOut_valid : std_logic;
  signal cond_br21_falseOut_ready : std_logic;
  signal buffer62_outs_valid : std_logic;
  signal buffer62_outs_ready : std_logic;
  signal buffer63_outs_valid : std_logic;
  signal buffer63_outs_ready : std_logic;
  signal buffer64_outs_valid : std_logic;
  signal buffer64_outs_ready : std_logic;
  signal buffer65_outs_valid : std_logic;
  signal buffer65_outs_ready : std_logic;
  signal buffer66_outs_valid : std_logic;
  signal buffer66_outs_ready : std_logic;
  signal buffer211_outs : std_logic_vector(0 downto 0);
  signal buffer211_outs_valid : std_logic;
  signal buffer211_outs_ready : std_logic;
  signal buffer212_outs : std_logic_vector(0 downto 0);
  signal buffer212_outs_valid : std_logic;
  signal buffer212_outs_ready : std_logic;
  signal buffer213_outs : std_logic_vector(0 downto 0);
  signal buffer213_outs_valid : std_logic;
  signal buffer213_outs_ready : std_logic;
  signal buffer214_outs : std_logic_vector(0 downto 0);
  signal buffer214_outs_valid : std_logic;
  signal buffer214_outs_ready : std_logic;
  signal buffer215_outs : std_logic_vector(0 downto 0);
  signal buffer215_outs_valid : std_logic;
  signal buffer215_outs_ready : std_logic;
  signal cond_br22_trueOut_valid : std_logic;
  signal cond_br22_trueOut_ready : std_logic;
  signal cond_br22_falseOut_valid : std_logic;
  signal cond_br22_falseOut_ready : std_logic;
  signal buffer5_outs_valid : std_logic;
  signal buffer5_outs_ready : std_logic;
  signal buffer6_outs_valid : std_logic;
  signal buffer6_outs_ready : std_logic;
  signal buffer7_outs_valid : std_logic;
  signal buffer7_outs_ready : std_logic;
  signal buffer8_outs_valid : std_logic;
  signal buffer8_outs_ready : std_logic;
  signal buffer9_outs_valid : std_logic;
  signal buffer9_outs_ready : std_logic;
  signal constant11_outs : std_logic_vector(1 downto 0);
  signal constant11_outs_valid : std_logic;
  signal constant11_outs_ready : std_logic;
  signal extsi4_outs : std_logic_vector(31 downto 0);
  signal extsi4_outs_valid : std_logic;
  signal extsi4_outs_ready : std_logic;
  signal buffer57_outs_valid : std_logic;
  signal buffer57_outs_ready : std_logic;
  signal buffer58_outs_valid : std_logic;
  signal buffer58_outs_ready : std_logic;
  signal buffer59_outs_valid : std_logic;
  signal buffer59_outs_ready : std_logic;
  signal buffer60_outs_valid : std_logic;
  signal buffer60_outs_ready : std_logic;
  signal buffer61_outs_valid : std_logic;
  signal buffer61_outs_ready : std_logic;
  signal constant13_outs : std_logic_vector(5 downto 0);
  signal constant13_outs_valid : std_logic;
  signal constant13_outs_ready : std_logic;
  signal extsi15_outs : std_logic_vector(6 downto 0);
  signal extsi15_outs_valid : std_logic;
  signal extsi15_outs_ready : std_logic;
  signal buffer52_outs_valid : std_logic;
  signal buffer52_outs_ready : std_logic;
  signal buffer53_outs_valid : std_logic;
  signal buffer53_outs_ready : std_logic;
  signal buffer54_outs_valid : std_logic;
  signal buffer54_outs_ready : std_logic;
  signal buffer55_outs_valid : std_logic;
  signal buffer55_outs_ready : std_logic;
  signal buffer56_outs_valid : std_logic;
  signal buffer56_outs_ready : std_logic;
  signal constant14_outs : std_logic_vector(1 downto 0);
  signal constant14_outs_valid : std_logic;
  signal constant14_outs_ready : std_logic;
  signal extsi16_outs : std_logic_vector(6 downto 0);
  signal extsi16_outs_valid : std_logic;
  signal extsi16_outs_ready : std_logic;
  signal buffer98_outs : std_logic_vector(31 downto 0);
  signal buffer98_outs_valid : std_logic;
  signal buffer98_outs_ready : std_logic;
  signal buffer99_outs : std_logic_vector(31 downto 0);
  signal buffer99_outs_valid : std_logic;
  signal buffer99_outs_ready : std_logic;
  signal buffer100_outs : std_logic_vector(31 downto 0);
  signal buffer100_outs_valid : std_logic;
  signal buffer100_outs_ready : std_logic;
  signal buffer101_outs : std_logic_vector(31 downto 0);
  signal buffer101_outs_valid : std_logic;
  signal buffer101_outs_ready : std_logic;
  signal buffer102_outs : std_logic_vector(31 downto 0);
  signal buffer102_outs_valid : std_logic;
  signal buffer102_outs_ready : std_logic;
  signal store0_addrOut : std_logic_vector(4 downto 0);
  signal store0_addrOut_valid : std_logic;
  signal store0_addrOut_ready : std_logic;
  signal store0_dataToMem : std_logic_vector(31 downto 0);
  signal store0_dataToMem_valid : std_logic;
  signal store0_dataToMem_ready : std_logic;
  signal addi2_result : std_logic_vector(6 downto 0);
  signal addi2_result_valid : std_logic;
  signal addi2_result_ready : std_logic;
  signal fork11_outs_0 : std_logic_vector(6 downto 0);
  signal fork11_outs_0_valid : std_logic;
  signal fork11_outs_0_ready : std_logic;
  signal fork11_outs_1 : std_logic_vector(6 downto 0);
  signal fork11_outs_1_valid : std_logic;
  signal fork11_outs_1_ready : std_logic;
  signal buffer191_outs : std_logic_vector(6 downto 0);
  signal buffer191_outs_valid : std_logic;
  signal buffer191_outs_ready : std_logic;
  signal buffer192_outs : std_logic_vector(6 downto 0);
  signal buffer192_outs_valid : std_logic;
  signal buffer192_outs_ready : std_logic;
  signal buffer193_outs : std_logic_vector(6 downto 0);
  signal buffer193_outs_valid : std_logic;
  signal buffer193_outs_ready : std_logic;
  signal buffer194_outs : std_logic_vector(6 downto 0);
  signal buffer194_outs_valid : std_logic;
  signal buffer194_outs_ready : std_logic;
  signal buffer195_outs : std_logic_vector(6 downto 0);
  signal buffer195_outs_valid : std_logic;
  signal buffer195_outs_ready : std_logic;
  signal trunci2_outs : std_logic_vector(5 downto 0);
  signal trunci2_outs_valid : std_logic;
  signal trunci2_outs_ready : std_logic;
  signal buffer186_outs : std_logic_vector(6 downto 0);
  signal buffer186_outs_valid : std_logic;
  signal buffer186_outs_ready : std_logic;
  signal buffer187_outs : std_logic_vector(6 downto 0);
  signal buffer187_outs_valid : std_logic;
  signal buffer187_outs_ready : std_logic;
  signal buffer188_outs : std_logic_vector(6 downto 0);
  signal buffer188_outs_valid : std_logic;
  signal buffer188_outs_ready : std_logic;
  signal buffer189_outs : std_logic_vector(6 downto 0);
  signal buffer189_outs_valid : std_logic;
  signal buffer189_outs_ready : std_logic;
  signal buffer190_outs : std_logic_vector(6 downto 0);
  signal buffer190_outs_valid : std_logic;
  signal buffer190_outs_ready : std_logic;
  signal cmpi1_result : std_logic_vector(0 downto 0);
  signal cmpi1_result_valid : std_logic;
  signal cmpi1_result_ready : std_logic;
  signal fork12_outs_0 : std_logic_vector(0 downto 0);
  signal fork12_outs_0_valid : std_logic;
  signal fork12_outs_0_ready : std_logic;
  signal fork12_outs_1 : std_logic_vector(0 downto 0);
  signal fork12_outs_1_valid : std_logic;
  signal fork12_outs_1_ready : std_logic;
  signal fork12_outs_2 : std_logic_vector(0 downto 0);
  signal fork12_outs_2_valid : std_logic;
  signal fork12_outs_2_ready : std_logic;
  signal fork12_outs_3 : std_logic_vector(0 downto 0);
  signal fork12_outs_3_valid : std_logic;
  signal fork12_outs_3_ready : std_logic;
  signal buffer0_outs_valid : std_logic;
  signal buffer0_outs_ready : std_logic;
  signal buffer1_outs_valid : std_logic;
  signal buffer1_outs_ready : std_logic;
  signal buffer2_outs_valid : std_logic;
  signal buffer2_outs_ready : std_logic;
  signal buffer3_outs_valid : std_logic;
  signal buffer3_outs_ready : std_logic;
  signal buffer4_outs_valid : std_logic;
  signal buffer4_outs_ready : std_logic;

begin

  out0 <= cond_br20_falseOut;
  out0_valid <= cond_br20_falseOut_valid;
  cond_br20_falseOut_ready <= out0_ready;
  q_end_valid <= mem_controller1_memEnd_valid;
  mem_controller1_memEnd_ready <= q_end_ready;
  end_valid <= buffer4_outs_valid;
  buffer4_outs_ready <= end_ready;
  q_loadEn <= mem_controller1_loadEn;
  q_loadAddr <= mem_controller1_loadAddr;
  q_storeEn <= mem_controller1_storeEn;
  q_storeAddr <= mem_controller1_storeAddr;
  q_storeData <= mem_controller1_storeData;

  fork0 : entity work.handshake_fork_0(arch)
    port map(
      ins_valid => start_valid,
      ins_ready => start_ready,
      clk => clk,
      rst => rst,
      outs_valid(0) => fork0_outs_0_valid,
      outs_valid(1) => fork0_outs_1_valid,
      outs_valid(2) => fork0_outs_2_valid,
      outs_valid(3) => fork0_outs_3_valid,
      outs_valid(4) => fork0_outs_4_valid,
      outs_ready(0) => fork0_outs_0_ready,
      outs_ready(1) => fork0_outs_1_ready,
      outs_ready(2) => fork0_outs_2_ready,
      outs_ready(3) => fork0_outs_3_ready,
      outs_ready(4) => fork0_outs_4_ready
    );

  buffer20 : entity work.handshake_buffer_0(arch)
    port map(
      ins_valid => fork0_outs_4_valid,
      ins_ready => fork0_outs_4_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer20_outs_valid,
      outs_ready => buffer20_outs_ready
    );

  buffer21 : entity work.handshake_buffer_0(arch)
    port map(
      ins_valid => buffer20_outs_valid,
      ins_ready => buffer20_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer21_outs_valid,
      outs_ready => buffer21_outs_ready
    );

  buffer22 : entity work.handshake_buffer_0(arch)
    port map(
      ins_valid => buffer21_outs_valid,
      ins_ready => buffer21_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer22_outs_valid,
      outs_ready => buffer22_outs_ready
    );

  buffer23 : entity work.handshake_buffer_0(arch)
    port map(
      ins_valid => buffer22_outs_valid,
      ins_ready => buffer22_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer23_outs_valid,
      outs_ready => buffer23_outs_ready
    );

  buffer24 : entity work.handshake_buffer_0(arch)
    port map(
      ins_valid => buffer23_outs_valid,
      ins_ready => buffer23_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer24_outs_valid,
      outs_ready => buffer24_outs_ready
    );

  mem_controller1 : entity work.handshake_mem_controller_0(arch)
    port map(
      loadData => q_loadData,
      memStart_valid => q_start_valid,
      memStart_ready => q_start_ready,
      ctrl(0) => extsi4_outs,
      ctrl_valid(0) => extsi4_outs_valid,
      ctrl_ready(0) => extsi4_outs_ready,
      stAddr(0) => store0_addrOut,
      stAddr_valid(0) => store0_addrOut_valid,
      stAddr_ready(0) => store0_addrOut_ready,
      stData(0) => store0_dataToMem,
      stData_valid(0) => store0_dataToMem_valid,
      stData_ready(0) => store0_dataToMem_ready,
      ctrlEnd_valid => buffer24_outs_valid,
      ctrlEnd_ready => buffer24_outs_ready,
      clk => clk,
      rst => rst,
      memEnd_valid => mem_controller1_memEnd_valid,
      memEnd_ready => mem_controller1_memEnd_ready,
      loadEn => mem_controller1_loadEn,
      loadAddr => mem_controller1_loadAddr,
      storeEn => mem_controller1_storeEn,
      storeAddr => mem_controller1_storeAddr,
      storeData => mem_controller1_storeData
    );

  buffer15 : entity work.handshake_buffer_0(arch)
    port map(
      ins_valid => fork0_outs_3_valid,
      ins_ready => fork0_outs_3_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer15_outs_valid,
      outs_ready => buffer15_outs_ready
    );

  buffer16 : entity work.handshake_buffer_0(arch)
    port map(
      ins_valid => buffer15_outs_valid,
      ins_ready => buffer15_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer16_outs_valid,
      outs_ready => buffer16_outs_ready
    );

  buffer17 : entity work.handshake_buffer_0(arch)
    port map(
      ins_valid => buffer16_outs_valid,
      ins_ready => buffer16_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer17_outs_valid,
      outs_ready => buffer17_outs_ready
    );

  buffer18 : entity work.handshake_buffer_0(arch)
    port map(
      ins_valid => buffer17_outs_valid,
      ins_ready => buffer17_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer18_outs_valid,
      outs_ready => buffer18_outs_ready
    );

  buffer19 : entity work.handshake_buffer_0(arch)
    port map(
      ins_valid => buffer18_outs_valid,
      ins_ready => buffer18_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer19_outs_valid,
      outs_ready => buffer19_outs_ready
    );

  constant0 : entity work.handshake_constant_0(arch)
    port map(
      ctrl_valid => buffer19_outs_valid,
      ctrl_ready => buffer19_outs_ready,
      clk => clk,
      rst => rst,
      outs => constant0_outs,
      outs_valid => constant0_outs_valid,
      outs_ready => constant0_outs_ready
    );

  fork1 : entity work.handshake_fork_1(arch)
    port map(
      ins => constant0_outs,
      ins_valid => constant0_outs_valid,
      ins_ready => constant0_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork1_outs_0,
      outs(1) => fork1_outs_1,
      outs_valid(0) => fork1_outs_0_valid,
      outs_valid(1) => fork1_outs_1_valid,
      outs_ready(0) => fork1_outs_0_ready,
      outs_ready(1) => fork1_outs_1_ready
    );

  buffer30 : entity work.handshake_buffer_1(arch)
    port map(
      ins => fork1_outs_1,
      ins_valid => fork1_outs_1_valid,
      ins_ready => fork1_outs_1_ready,
      clk => clk,
      rst => rst,
      outs => buffer30_outs,
      outs_valid => buffer30_outs_valid,
      outs_ready => buffer30_outs_ready
    );

  buffer31 : entity work.handshake_buffer_1(arch)
    port map(
      ins => buffer30_outs,
      ins_valid => buffer30_outs_valid,
      ins_ready => buffer30_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer31_outs,
      outs_valid => buffer31_outs_valid,
      outs_ready => buffer31_outs_ready
    );

  buffer32 : entity work.handshake_buffer_1(arch)
    port map(
      ins => buffer31_outs,
      ins_valid => buffer31_outs_valid,
      ins_ready => buffer31_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer32_outs,
      outs_valid => buffer32_outs_valid,
      outs_ready => buffer32_outs_ready
    );

  buffer33 : entity work.handshake_buffer_1(arch)
    port map(
      ins => buffer32_outs,
      ins_valid => buffer32_outs_valid,
      ins_ready => buffer32_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer33_outs,
      outs_valid => buffer33_outs_valid,
      outs_ready => buffer33_outs_ready
    );

  buffer34 : entity work.handshake_buffer_1(arch)
    port map(
      ins => buffer33_outs,
      ins_valid => buffer33_outs_valid,
      ins_ready => buffer33_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer34_outs,
      outs_valid => buffer34_outs_valid,
      outs_ready => buffer34_outs_ready
    );

  extsi7 : entity work.handshake_extsi_0(arch)
    port map(
      ins => buffer34_outs,
      ins_valid => buffer34_outs_valid,
      ins_ready => buffer34_outs_ready,
      clk => clk,
      rst => rst,
      outs => extsi7_outs,
      outs_valid => extsi7_outs_valid,
      outs_ready => extsi7_outs_ready
    );

  buffer25 : entity work.handshake_buffer_1(arch)
    port map(
      ins => fork1_outs_0,
      ins_valid => fork1_outs_0_valid,
      ins_ready => fork1_outs_0_ready,
      clk => clk,
      rst => rst,
      outs => buffer25_outs,
      outs_valid => buffer25_outs_valid,
      outs_ready => buffer25_outs_ready
    );

  buffer26 : entity work.handshake_buffer_1(arch)
    port map(
      ins => buffer25_outs,
      ins_valid => buffer25_outs_valid,
      ins_ready => buffer25_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer26_outs,
      outs_valid => buffer26_outs_valid,
      outs_ready => buffer26_outs_ready
    );

  buffer27 : entity work.handshake_buffer_1(arch)
    port map(
      ins => buffer26_outs,
      ins_valid => buffer26_outs_valid,
      ins_ready => buffer26_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer27_outs,
      outs_valid => buffer27_outs_valid,
      outs_ready => buffer27_outs_ready
    );

  buffer28 : entity work.handshake_buffer_1(arch)
    port map(
      ins => buffer27_outs,
      ins_valid => buffer27_outs_valid,
      ins_ready => buffer27_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer28_outs,
      outs_valid => buffer28_outs_valid,
      outs_ready => buffer28_outs_ready
    );

  buffer29 : entity work.handshake_buffer_1(arch)
    port map(
      ins => buffer28_outs,
      ins_valid => buffer28_outs_valid,
      ins_ready => buffer28_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer29_outs,
      outs_valid => buffer29_outs_valid,
      outs_ready => buffer29_outs_ready
    );

  buffer196 : entity work.handshake_buffer_1(arch)
    port map(
      ins => fork12_outs_0,
      ins_valid => fork12_outs_0_valid,
      ins_ready => fork12_outs_0_ready,
      clk => clk,
      rst => rst,
      outs => buffer196_outs,
      outs_valid => buffer196_outs_valid,
      outs_ready => buffer196_outs_ready
    );

  buffer197 : entity work.handshake_buffer_1(arch)
    port map(
      ins => buffer196_outs,
      ins_valid => buffer196_outs_valid,
      ins_ready => buffer196_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer197_outs,
      outs_valid => buffer197_outs_valid,
      outs_ready => buffer197_outs_ready
    );

  buffer198 : entity work.handshake_buffer_1(arch)
    port map(
      ins => buffer197_outs,
      ins_valid => buffer197_outs_valid,
      ins_ready => buffer197_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer198_outs,
      outs_valid => buffer198_outs_valid,
      outs_ready => buffer198_outs_ready
    );

  buffer199 : entity work.handshake_buffer_1(arch)
    port map(
      ins => buffer198_outs,
      ins_valid => buffer198_outs_valid,
      ins_ready => buffer198_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer199_outs,
      outs_valid => buffer199_outs_valid,
      outs_ready => buffer199_outs_ready
    );

  buffer200 : entity work.handshake_buffer_1(arch)
    port map(
      ins => buffer199_outs,
      ins_valid => buffer199_outs_valid,
      ins_ready => buffer199_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer200_outs,
      outs_valid => buffer200_outs_valid,
      outs_ready => buffer200_outs_ready
    );

  merge0 : entity work.handshake_merge_0(arch)
    port map(
      ins(0) => buffer29_outs,
      ins(1) => buffer200_outs,
      ins_valid(0) => buffer29_outs_valid,
      ins_valid(1) => buffer200_outs_valid,
      ins_ready(0) => buffer29_outs_ready,
      ins_ready(1) => buffer200_outs_ready,
      clk => clk,
      rst => rst,
      outs => merge0_outs,
      outs_valid => merge0_outs_valid,
      outs_ready => merge0_outs_ready
    );

  buffer35 : entity work.handshake_buffer_1(arch)
    port map(
      ins => merge0_outs,
      ins_valid => merge0_outs_valid,
      ins_ready => merge0_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer35_outs,
      outs_valid => buffer35_outs_valid,
      outs_ready => buffer35_outs_ready
    );

  fork2 : entity work.handshake_fork_1(arch)
    port map(
      ins => buffer35_outs,
      ins_valid => buffer35_outs_valid,
      ins_ready => buffer35_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork2_outs_0,
      outs(1) => fork2_outs_1,
      outs_valid(0) => fork2_outs_0_valid,
      outs_valid(1) => fork2_outs_1_valid,
      outs_ready(0) => fork2_outs_0_ready,
      outs_ready(1) => fork2_outs_1_ready
    );

  buffer10 : entity work.handshake_buffer_0(arch)
    port map(
      ins_valid => fork0_outs_2_valid,
      ins_ready => fork0_outs_2_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer10_outs_valid,
      outs_ready => buffer10_outs_ready
    );

  buffer11 : entity work.handshake_buffer_0(arch)
    port map(
      ins_valid => buffer10_outs_valid,
      ins_ready => buffer10_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer11_outs_valid,
      outs_ready => buffer11_outs_ready
    );

  buffer12 : entity work.handshake_buffer_0(arch)
    port map(
      ins_valid => buffer11_outs_valid,
      ins_ready => buffer11_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer12_outs_valid,
      outs_ready => buffer12_outs_ready
    );

  buffer13 : entity work.handshake_buffer_0(arch)
    port map(
      ins_valid => buffer12_outs_valid,
      ins_ready => buffer12_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer13_outs_valid,
      outs_ready => buffer13_outs_ready
    );

  buffer14 : entity work.handshake_buffer_0(arch)
    port map(
      ins_valid => buffer13_outs_valid,
      ins_ready => buffer13_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer14_outs_valid,
      outs_ready => buffer14_outs_ready
    );

  buffer41 : entity work.handshake_buffer_1(arch)
    port map(
      ins => fork2_outs_1,
      ins_valid => fork2_outs_1_valid,
      ins_ready => fork2_outs_1_ready,
      clk => clk,
      rst => rst,
      outs => buffer41_outs,
      outs_valid => buffer41_outs_valid,
      outs_ready => buffer41_outs_ready
    );

  buffer42 : entity work.handshake_buffer_1(arch)
    port map(
      ins => buffer41_outs,
      ins_valid => buffer41_outs_valid,
      ins_ready => buffer41_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer42_outs,
      outs_valid => buffer42_outs_valid,
      outs_ready => buffer42_outs_ready
    );

  buffer43 : entity work.handshake_buffer_1(arch)
    port map(
      ins => buffer42_outs,
      ins_valid => buffer42_outs_valid,
      ins_ready => buffer42_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer43_outs,
      outs_valid => buffer43_outs_valid,
      outs_ready => buffer43_outs_ready
    );

  buffer44 : entity work.handshake_buffer_1(arch)
    port map(
      ins => buffer43_outs,
      ins_valid => buffer43_outs_valid,
      ins_ready => buffer43_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer44_outs,
      outs_valid => buffer44_outs_valid,
      outs_ready => buffer44_outs_ready
    );

  buffer45 : entity work.handshake_buffer_1(arch)
    port map(
      ins => buffer44_outs,
      ins_valid => buffer44_outs_valid,
      ins_ready => buffer44_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer45_outs,
      outs_valid => buffer45_outs_valid,
      outs_ready => buffer45_outs_ready
    );

  mux0 : entity work.handshake_mux_0(arch)
    port map(
      index => buffer45_outs,
      index_valid => buffer45_outs_valid,
      index_ready => buffer45_outs_ready,
      ins_valid(0) => buffer14_outs_valid,
      ins_valid(1) => cond_br22_trueOut_valid,
      ins_ready(0) => buffer14_outs_ready,
      ins_ready(1) => cond_br22_trueOut_ready,
      clk => clk,
      rst => rst,
      outs_valid => mux0_outs_valid,
      outs_ready => mux0_outs_ready
    );

  buffer46 : entity work.handshake_buffer_2(arch)
    port map(
      ins_valid => mux0_outs_valid,
      ins_ready => mux0_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer46_outs_valid,
      outs_ready => buffer46_outs_ready
    );

  buffer47 : entity work.handshake_buffer_0(arch)
    port map(
      ins_valid => buffer46_outs_valid,
      ins_ready => buffer46_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer47_outs_valid,
      outs_ready => buffer47_outs_ready
    );

  buffer48 : entity work.handshake_buffer_0(arch)
    port map(
      ins_valid => buffer47_outs_valid,
      ins_ready => buffer47_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer48_outs_valid,
      outs_ready => buffer48_outs_ready
    );

  buffer49 : entity work.handshake_buffer_0(arch)
    port map(
      ins_valid => buffer48_outs_valid,
      ins_ready => buffer48_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer49_outs_valid,
      outs_ready => buffer49_outs_ready
    );

  buffer50 : entity work.handshake_buffer_0(arch)
    port map(
      ins_valid => buffer49_outs_valid,
      ins_ready => buffer49_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer50_outs_valid,
      outs_ready => buffer50_outs_ready
    );

  buffer51 : entity work.handshake_buffer_0(arch)
    port map(
      ins_valid => buffer50_outs_valid,
      ins_ready => buffer50_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer51_outs_valid,
      outs_ready => buffer51_outs_ready
    );

  fork3 : entity work.handshake_fork_0(arch)
    port map(
      ins_valid => buffer51_outs_valid,
      ins_ready => buffer51_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid(0) => fork3_outs_0_valid,
      outs_valid(1) => fork3_outs_1_valid,
      outs_valid(2) => fork3_outs_2_valid,
      outs_valid(3) => fork3_outs_3_valid,
      outs_valid(4) => fork3_outs_4_valid,
      outs_ready(0) => fork3_outs_0_ready,
      outs_ready(1) => fork3_outs_1_ready,
      outs_ready(2) => fork3_outs_2_ready,
      outs_ready(3) => fork3_outs_3_ready,
      outs_ready(4) => fork3_outs_4_ready
    );

  buffer36 : entity work.handshake_buffer_1(arch)
    port map(
      ins => fork2_outs_0,
      ins_valid => fork2_outs_0_valid,
      ins_ready => fork2_outs_0_ready,
      clk => clk,
      rst => rst,
      outs => buffer36_outs,
      outs_valid => buffer36_outs_valid,
      outs_ready => buffer36_outs_ready
    );

  buffer37 : entity work.handshake_buffer_1(arch)
    port map(
      ins => buffer36_outs,
      ins_valid => buffer36_outs_valid,
      ins_ready => buffer36_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer37_outs,
      outs_valid => buffer37_outs_valid,
      outs_ready => buffer37_outs_ready
    );

  buffer38 : entity work.handshake_buffer_1(arch)
    port map(
      ins => buffer37_outs,
      ins_valid => buffer37_outs_valid,
      ins_ready => buffer37_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer38_outs,
      outs_valid => buffer38_outs_valid,
      outs_ready => buffer38_outs_ready
    );

  buffer39 : entity work.handshake_buffer_1(arch)
    port map(
      ins => buffer38_outs,
      ins_valid => buffer38_outs_valid,
      ins_ready => buffer38_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer39_outs,
      outs_valid => buffer39_outs_valid,
      outs_ready => buffer39_outs_ready
    );

  buffer40 : entity work.handshake_buffer_1(arch)
    port map(
      ins => buffer39_outs,
      ins_valid => buffer39_outs_valid,
      ins_ready => buffer39_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer40_outs,
      outs_valid => buffer40_outs_valid,
      outs_ready => buffer40_outs_ready
    );

  mux5 : entity work.handshake_mux_1(arch)
    port map(
      index => buffer40_outs,
      index_valid => buffer40_outs_valid,
      index_ready => buffer40_outs_ready,
      ins(0) => extsi7_outs,
      ins(1) => cond_br21_trueOut,
      ins_valid(0) => extsi7_outs_valid,
      ins_valid(1) => cond_br21_trueOut_valid,
      ins_ready(0) => extsi7_outs_ready,
      ins_ready(1) => cond_br21_trueOut_ready,
      clk => clk,
      rst => rst,
      outs => mux5_outs,
      outs_valid => mux5_outs_valid,
      outs_ready => mux5_outs_ready
    );

  buffer77 : entity work.handshake_buffer_3(arch)
    port map(
      ins => mux5_outs,
      ins_valid => mux5_outs_valid,
      ins_ready => mux5_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer77_outs,
      outs_valid => buffer77_outs_valid,
      outs_ready => buffer77_outs_ready
    );

  buffer78 : entity work.handshake_buffer_4(arch)
    port map(
      ins => buffer77_outs,
      ins_valid => buffer77_outs_valid,
      ins_ready => buffer77_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer78_outs,
      outs_valid => buffer78_outs_valid,
      outs_ready => buffer78_outs_ready
    );

  buffer79 : entity work.handshake_buffer_4(arch)
    port map(
      ins => buffer78_outs,
      ins_valid => buffer78_outs_valid,
      ins_ready => buffer78_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer79_outs,
      outs_valid => buffer79_outs_valid,
      outs_ready => buffer79_outs_ready
    );

  buffer80 : entity work.handshake_buffer_4(arch)
    port map(
      ins => buffer79_outs,
      ins_valid => buffer79_outs_valid,
      ins_ready => buffer79_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer80_outs,
      outs_valid => buffer80_outs_valid,
      outs_ready => buffer80_outs_ready
    );

  buffer81 : entity work.handshake_buffer_4(arch)
    port map(
      ins => buffer80_outs,
      ins_valid => buffer80_outs_valid,
      ins_ready => buffer80_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer81_outs,
      outs_valid => buffer81_outs_valid,
      outs_ready => buffer81_outs_ready
    );

  buffer82 : entity work.handshake_buffer_4(arch)
    port map(
      ins => buffer81_outs,
      ins_valid => buffer81_outs_valid,
      ins_ready => buffer81_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer82_outs,
      outs_valid => buffer82_outs_valid,
      outs_ready => buffer82_outs_ready
    );

  fork4 : entity work.handshake_fork_2(arch)
    port map(
      ins => buffer82_outs,
      ins_valid => buffer82_outs_valid,
      ins_ready => buffer82_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork4_outs_0,
      outs(1) => fork4_outs_1,
      outs(2) => fork4_outs_2,
      outs_valid(0) => fork4_outs_0_valid,
      outs_valid(1) => fork4_outs_1_valid,
      outs_valid(2) => fork4_outs_2_valid,
      outs_ready(0) => fork4_outs_0_ready,
      outs_ready(1) => fork4_outs_1_ready,
      outs_ready(2) => fork4_outs_2_ready
    );

  buffer93 : entity work.handshake_buffer_4(arch)
    port map(
      ins => fork4_outs_2,
      ins_valid => fork4_outs_2_valid,
      ins_ready => fork4_outs_2_ready,
      clk => clk,
      rst => rst,
      outs => buffer93_outs,
      outs_valid => buffer93_outs_valid,
      outs_ready => buffer93_outs_ready
    );

  buffer94 : entity work.handshake_buffer_4(arch)
    port map(
      ins => buffer93_outs,
      ins_valid => buffer93_outs_valid,
      ins_ready => buffer93_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer94_outs,
      outs_valid => buffer94_outs_valid,
      outs_ready => buffer94_outs_ready
    );

  buffer95 : entity work.handshake_buffer_4(arch)
    port map(
      ins => buffer94_outs,
      ins_valid => buffer94_outs_valid,
      ins_ready => buffer94_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer95_outs,
      outs_valid => buffer95_outs_valid,
      outs_ready => buffer95_outs_ready
    );

  buffer96 : entity work.handshake_buffer_4(arch)
    port map(
      ins => buffer95_outs,
      ins_valid => buffer95_outs_valid,
      ins_ready => buffer95_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer96_outs,
      outs_valid => buffer96_outs_valid,
      outs_ready => buffer96_outs_ready
    );

  buffer97 : entity work.handshake_buffer_4(arch)
    port map(
      ins => buffer96_outs,
      ins_valid => buffer96_outs_valid,
      ins_ready => buffer96_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer97_outs,
      outs_valid => buffer97_outs_valid,
      outs_ready => buffer97_outs_ready
    );

  extsi8 : entity work.handshake_extsi_1(arch)
    port map(
      ins => buffer97_outs,
      ins_valid => buffer97_outs_valid,
      ins_ready => buffer97_outs_ready,
      clk => clk,
      rst => rst,
      outs => extsi8_outs,
      outs_valid => extsi8_outs_valid,
      outs_ready => extsi8_outs_ready
    );

  buffer88 : entity work.handshake_buffer_4(arch)
    port map(
      ins => fork4_outs_1,
      ins_valid => fork4_outs_1_valid,
      ins_ready => fork4_outs_1_ready,
      clk => clk,
      rst => rst,
      outs => buffer88_outs,
      outs_valid => buffer88_outs_valid,
      outs_ready => buffer88_outs_ready
    );

  buffer89 : entity work.handshake_buffer_4(arch)
    port map(
      ins => buffer88_outs,
      ins_valid => buffer88_outs_valid,
      ins_ready => buffer88_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer89_outs,
      outs_valid => buffer89_outs_valid,
      outs_ready => buffer89_outs_ready
    );

  buffer90 : entity work.handshake_buffer_4(arch)
    port map(
      ins => buffer89_outs,
      ins_valid => buffer89_outs_valid,
      ins_ready => buffer89_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer90_outs,
      outs_valid => buffer90_outs_valid,
      outs_ready => buffer90_outs_ready
    );

  buffer91 : entity work.handshake_buffer_4(arch)
    port map(
      ins => buffer90_outs,
      ins_valid => buffer90_outs_valid,
      ins_ready => buffer90_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer91_outs,
      outs_valid => buffer91_outs_valid,
      outs_ready => buffer91_outs_ready
    );

  buffer92 : entity work.handshake_buffer_4(arch)
    port map(
      ins => buffer91_outs,
      ins_valid => buffer91_outs_valid,
      ins_ready => buffer91_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer92_outs,
      outs_valid => buffer92_outs_valid,
      outs_ready => buffer92_outs_ready
    );

  extsi9 : entity work.handshake_extsi_2(arch)
    port map(
      ins => buffer92_outs,
      ins_valid => buffer92_outs_valid,
      ins_ready => buffer92_outs_ready,
      clk => clk,
      rst => rst,
      outs => extsi9_outs,
      outs_valid => extsi9_outs_valid,
      outs_ready => extsi9_outs_ready
    );

  buffer83 : entity work.handshake_buffer_4(arch)
    port map(
      ins => fork4_outs_0,
      ins_valid => fork4_outs_0_valid,
      ins_ready => fork4_outs_0_ready,
      clk => clk,
      rst => rst,
      outs => buffer83_outs,
      outs_valid => buffer83_outs_valid,
      outs_ready => buffer83_outs_ready
    );

  buffer84 : entity work.handshake_buffer_4(arch)
    port map(
      ins => buffer83_outs,
      ins_valid => buffer83_outs_valid,
      ins_ready => buffer83_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer84_outs,
      outs_valid => buffer84_outs_valid,
      outs_ready => buffer84_outs_ready
    );

  buffer85 : entity work.handshake_buffer_4(arch)
    port map(
      ins => buffer84_outs,
      ins_valid => buffer84_outs_valid,
      ins_ready => buffer84_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer85_outs,
      outs_valid => buffer85_outs_valid,
      outs_ready => buffer85_outs_ready
    );

  buffer86 : entity work.handshake_buffer_4(arch)
    port map(
      ins => buffer85_outs,
      ins_valid => buffer85_outs_valid,
      ins_ready => buffer85_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer86_outs,
      outs_valid => buffer86_outs_valid,
      outs_ready => buffer86_outs_ready
    );

  buffer87 : entity work.handshake_buffer_4(arch)
    port map(
      ins => buffer86_outs,
      ins_valid => buffer86_outs_valid,
      ins_ready => buffer86_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer87_outs,
      outs_valid => buffer87_outs_valid,
      outs_ready => buffer87_outs_ready
    );

  trunci0 : entity work.handshake_trunci_0(arch)
    port map(
      ins => buffer87_outs,
      ins_valid => buffer87_outs_valid,
      ins_ready => buffer87_outs_ready,
      clk => clk,
      rst => rst,
      outs => trunci0_outs,
      outs_valid => trunci0_outs_valid,
      outs_ready => trunci0_outs_ready
    );

  buffer72 : entity work.handshake_buffer_0(arch)
    port map(
      ins_valid => fork3_outs_4_valid,
      ins_ready => fork3_outs_4_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer72_outs_valid,
      outs_ready => buffer72_outs_ready
    );

  buffer73 : entity work.handshake_buffer_0(arch)
    port map(
      ins_valid => buffer72_outs_valid,
      ins_ready => buffer72_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer73_outs_valid,
      outs_ready => buffer73_outs_ready
    );

  buffer74 : entity work.handshake_buffer_0(arch)
    port map(
      ins_valid => buffer73_outs_valid,
      ins_ready => buffer73_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer74_outs_valid,
      outs_ready => buffer74_outs_ready
    );

  buffer75 : entity work.handshake_buffer_0(arch)
    port map(
      ins_valid => buffer74_outs_valid,
      ins_ready => buffer74_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer75_outs_valid,
      outs_ready => buffer75_outs_ready
    );

  buffer76 : entity work.handshake_buffer_0(arch)
    port map(
      ins_valid => buffer75_outs_valid,
      ins_ready => buffer75_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer76_outs_valid,
      outs_ready => buffer76_outs_ready
    );

  constant8 : entity work.handshake_constant_0(arch)
    port map(
      ctrl_valid => buffer76_outs_valid,
      ctrl_ready => buffer76_outs_ready,
      clk => clk,
      rst => rst,
      outs => constant8_outs,
      outs_valid => constant8_outs_valid,
      outs_ready => constant8_outs_ready
    );

  extsi10 : entity work.handshake_extsi_0(arch)
    port map(
      ins => constant8_outs,
      ins_valid => constant8_outs_valid,
      ins_ready => constant8_outs_ready,
      clk => clk,
      rst => rst,
      outs => extsi10_outs,
      outs_valid => extsi10_outs_valid,
      outs_ready => extsi10_outs_ready
    );

  buffer171 : entity work.handshake_buffer_1(arch)
    port map(
      ins => fork10_outs_0,
      ins_valid => fork10_outs_0_valid,
      ins_ready => fork10_outs_0_ready,
      clk => clk,
      rst => rst,
      outs => buffer171_outs,
      outs_valid => buffer171_outs_valid,
      outs_ready => buffer171_outs_ready
    );

  buffer172 : entity work.handshake_buffer_1(arch)
    port map(
      ins => buffer171_outs,
      ins_valid => buffer171_outs_valid,
      ins_ready => buffer171_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer172_outs,
      outs_valid => buffer172_outs_valid,
      outs_ready => buffer172_outs_ready
    );

  buffer173 : entity work.handshake_buffer_1(arch)
    port map(
      ins => buffer172_outs,
      ins_valid => buffer172_outs_valid,
      ins_ready => buffer172_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer173_outs,
      outs_valid => buffer173_outs_valid,
      outs_ready => buffer173_outs_ready
    );

  buffer174 : entity work.handshake_buffer_1(arch)
    port map(
      ins => buffer173_outs,
      ins_valid => buffer173_outs_valid,
      ins_ready => buffer173_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer174_outs,
      outs_valid => buffer174_outs_valid,
      outs_ready => buffer174_outs_ready
    );

  buffer175 : entity work.handshake_buffer_1(arch)
    port map(
      ins => buffer174_outs,
      ins_valid => buffer174_outs_valid,
      ins_ready => buffer174_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer175_outs,
      outs_valid => buffer175_outs_valid,
      outs_ready => buffer175_outs_ready
    );

  cond_br17 : entity work.handshake_cond_br_0(arch)
    port map(
      condition => buffer175_outs,
      condition_valid => buffer175_outs_valid,
      condition_ready => buffer175_outs_ready,
      data => muli0_result,
      data_valid => muli0_result_valid,
      data_ready => muli0_result_ready,
      clk => clk,
      rst => rst,
      trueOut => cond_br17_trueOut,
      trueOut_valid => cond_br17_trueOut_valid,
      trueOut_ready => cond_br17_trueOut_ready,
      falseOut => cond_br17_falseOut,
      falseOut_valid => cond_br17_falseOut_valid,
      falseOut_ready => cond_br17_falseOut_ready
    );

  fork5 : entity work.handshake_fork_3(arch)
    port map(
      ins => cond_br17_falseOut,
      ins_valid => cond_br17_falseOut_valid,
      ins_ready => cond_br17_falseOut_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork5_outs_0,
      outs(1) => fork5_outs_1,
      outs_valid(0) => fork5_outs_0_valid,
      outs_valid(1) => fork5_outs_1_valid,
      outs_ready(0) => fork5_outs_0_ready,
      outs_ready(1) => fork5_outs_1_ready
    );

  buffer176 : entity work.handshake_buffer_1(arch)
    port map(
      ins => fork10_outs_1,
      ins_valid => fork10_outs_1_valid,
      ins_ready => fork10_outs_1_ready,
      clk => clk,
      rst => rst,
      outs => buffer176_outs,
      outs_valid => buffer176_outs_valid,
      outs_ready => buffer176_outs_ready
    );

  buffer177 : entity work.handshake_buffer_1(arch)
    port map(
      ins => buffer176_outs,
      ins_valid => buffer176_outs_valid,
      ins_ready => buffer176_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer177_outs,
      outs_valid => buffer177_outs_valid,
      outs_ready => buffer177_outs_ready
    );

  buffer178 : entity work.handshake_buffer_1(arch)
    port map(
      ins => buffer177_outs,
      ins_valid => buffer177_outs_valid,
      ins_ready => buffer177_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer178_outs,
      outs_valid => buffer178_outs_valid,
      outs_ready => buffer178_outs_ready
    );

  buffer179 : entity work.handshake_buffer_1(arch)
    port map(
      ins => buffer178_outs,
      ins_valid => buffer178_outs_valid,
      ins_ready => buffer178_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer179_outs,
      outs_valid => buffer179_outs_valid,
      outs_ready => buffer179_outs_ready
    );

  buffer180 : entity work.handshake_buffer_1(arch)
    port map(
      ins => buffer179_outs,
      ins_valid => buffer179_outs_valid,
      ins_ready => buffer179_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer180_outs,
      outs_valid => buffer180_outs_valid,
      outs_ready => buffer180_outs_ready
    );

  cond_br18 : entity work.handshake_cond_br_1(arch)
    port map(
      condition => buffer180_outs,
      condition_valid => buffer180_outs_valid,
      condition_ready => buffer180_outs_ready,
      data => trunci1_outs,
      data_valid => trunci1_outs_valid,
      data_ready => trunci1_outs_ready,
      clk => clk,
      rst => rst,
      trueOut => cond_br18_trueOut,
      trueOut_valid => cond_br18_trueOut_valid,
      trueOut_ready => cond_br18_trueOut_ready,
      falseOut => cond_br18_falseOut,
      falseOut_valid => cond_br18_falseOut_valid,
      falseOut_ready => cond_br18_falseOut_ready
    );

  sink0 : entity work.handshake_sink_0(arch)
    port map(
      ins => cond_br18_falseOut,
      ins_valid => cond_br18_falseOut_valid,
      ins_ready => cond_br18_falseOut_ready,
      clk => clk,
      rst => rst
    );

  buffer134 : entity work.handshake_buffer_0(arch)
    port map(
      ins_valid => fork7_outs_2_valid,
      ins_ready => fork7_outs_2_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer134_outs_valid,
      outs_ready => buffer134_outs_ready
    );

  buffer135 : entity work.handshake_buffer_0(arch)
    port map(
      ins_valid => buffer134_outs_valid,
      ins_ready => buffer134_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer135_outs_valid,
      outs_ready => buffer135_outs_ready
    );

  buffer136 : entity work.handshake_buffer_0(arch)
    port map(
      ins_valid => buffer135_outs_valid,
      ins_ready => buffer135_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer136_outs_valid,
      outs_ready => buffer136_outs_ready
    );

  buffer137 : entity work.handshake_buffer_0(arch)
    port map(
      ins_valid => buffer136_outs_valid,
      ins_ready => buffer136_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer137_outs_valid,
      outs_ready => buffer137_outs_ready
    );

  buffer138 : entity work.handshake_buffer_0(arch)
    port map(
      ins_valid => buffer137_outs_valid,
      ins_ready => buffer137_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer138_outs_valid,
      outs_ready => buffer138_outs_ready
    );

  buffer181 : entity work.handshake_buffer_1(arch)
    port map(
      ins => fork10_outs_2,
      ins_valid => fork10_outs_2_valid,
      ins_ready => fork10_outs_2_ready,
      clk => clk,
      rst => rst,
      outs => buffer181_outs,
      outs_valid => buffer181_outs_valid,
      outs_ready => buffer181_outs_ready
    );

  buffer182 : entity work.handshake_buffer_1(arch)
    port map(
      ins => buffer181_outs,
      ins_valid => buffer181_outs_valid,
      ins_ready => buffer181_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer182_outs,
      outs_valid => buffer182_outs_valid,
      outs_ready => buffer182_outs_ready
    );

  buffer183 : entity work.handshake_buffer_1(arch)
    port map(
      ins => buffer182_outs,
      ins_valid => buffer182_outs_valid,
      ins_ready => buffer182_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer183_outs,
      outs_valid => buffer183_outs_valid,
      outs_ready => buffer183_outs_ready
    );

  buffer184 : entity work.handshake_buffer_1(arch)
    port map(
      ins => buffer183_outs,
      ins_valid => buffer183_outs_valid,
      ins_ready => buffer183_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer184_outs,
      outs_valid => buffer184_outs_valid,
      outs_ready => buffer184_outs_ready
    );

  buffer185 : entity work.handshake_buffer_1(arch)
    port map(
      ins => buffer184_outs,
      ins_valid => buffer184_outs_valid,
      ins_ready => buffer184_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer185_outs,
      outs_valid => buffer185_outs_valid,
      outs_ready => buffer185_outs_ready
    );

  cond_br19 : entity work.handshake_cond_br_2(arch)
    port map(
      condition => buffer185_outs,
      condition_valid => buffer185_outs_valid,
      condition_ready => buffer185_outs_ready,
      data_valid => buffer138_outs_valid,
      data_ready => buffer138_outs_ready,
      clk => clk,
      rst => rst,
      trueOut_valid => cond_br19_trueOut_valid,
      trueOut_ready => cond_br19_trueOut_ready,
      falseOut_valid => cond_br19_falseOut_valid,
      falseOut_ready => cond_br19_falseOut_ready
    );

  sink1 : entity work.handshake_sink_1(arch)
    port map(
      ins_valid => cond_br19_falseOut_valid,
      ins_ready => cond_br19_falseOut_ready,
      clk => clk,
      rst => rst
    );

  buffer67 : entity work.handshake_buffer_0(arch)
    port map(
      ins_valid => fork3_outs_3_valid,
      ins_ready => fork3_outs_3_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer67_outs_valid,
      outs_ready => buffer67_outs_ready
    );

  buffer68 : entity work.handshake_buffer_0(arch)
    port map(
      ins_valid => buffer67_outs_valid,
      ins_ready => buffer67_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer68_outs_valid,
      outs_ready => buffer68_outs_ready
    );

  buffer69 : entity work.handshake_buffer_0(arch)
    port map(
      ins_valid => buffer68_outs_valid,
      ins_ready => buffer68_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer69_outs_valid,
      outs_ready => buffer69_outs_ready
    );

  buffer70 : entity work.handshake_buffer_0(arch)
    port map(
      ins_valid => buffer69_outs_valid,
      ins_ready => buffer69_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer70_outs_valid,
      outs_ready => buffer70_outs_ready
    );

  buffer71 : entity work.handshake_buffer_0(arch)
    port map(
      ins_valid => buffer70_outs_valid,
      ins_ready => buffer70_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer71_outs_valid,
      outs_ready => buffer71_outs_ready
    );

  control_merge0 : entity work.handshake_control_merge_0(arch)
    port map(
      ins_valid(0) => buffer71_outs_valid,
      ins_valid(1) => cond_br19_trueOut_valid,
      ins_ready(0) => buffer71_outs_ready,
      ins_ready(1) => cond_br19_trueOut_ready,
      clk => clk,
      rst => rst,
      outs_valid => control_merge0_outs_valid,
      outs_ready => control_merge0_outs_ready,
      index => control_merge0_index,
      index_valid => control_merge0_index_valid,
      index_ready => control_merge0_index_ready
    );

  fork6 : entity work.handshake_fork_1(arch)
    port map(
      ins => control_merge0_index,
      ins_valid => control_merge0_index_valid,
      ins_ready => control_merge0_index_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork6_outs_0,
      outs(1) => fork6_outs_1,
      outs_valid(0) => fork6_outs_0_valid,
      outs_valid(1) => fork6_outs_1_valid,
      outs_ready(0) => fork6_outs_0_ready,
      outs_ready(1) => fork6_outs_1_ready
    );

  buffer108 : entity work.handshake_buffer_2(arch)
    port map(
      ins_valid => control_merge0_outs_valid,
      ins_ready => control_merge0_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer108_outs_valid,
      outs_ready => buffer108_outs_ready
    );

  buffer109 : entity work.handshake_buffer_0(arch)
    port map(
      ins_valid => buffer108_outs_valid,
      ins_ready => buffer108_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer109_outs_valid,
      outs_ready => buffer109_outs_ready
    );

  buffer110 : entity work.handshake_buffer_0(arch)
    port map(
      ins_valid => buffer109_outs_valid,
      ins_ready => buffer109_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer110_outs_valid,
      outs_ready => buffer110_outs_ready
    );

  buffer111 : entity work.handshake_buffer_0(arch)
    port map(
      ins_valid => buffer110_outs_valid,
      ins_ready => buffer110_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer111_outs_valid,
      outs_ready => buffer111_outs_ready
    );

  buffer112 : entity work.handshake_buffer_0(arch)
    port map(
      ins_valid => buffer111_outs_valid,
      ins_ready => buffer111_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer112_outs_valid,
      outs_ready => buffer112_outs_ready
    );

  buffer113 : entity work.handshake_buffer_0(arch)
    port map(
      ins_valid => buffer112_outs_valid,
      ins_ready => buffer112_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer113_outs_valid,
      outs_ready => buffer113_outs_ready
    );

  fork7 : entity work.handshake_fork_4(arch)
    port map(
      ins_valid => buffer113_outs_valid,
      ins_ready => buffer113_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid(0) => fork7_outs_0_valid,
      outs_valid(1) => fork7_outs_1_valid,
      outs_valid(2) => fork7_outs_2_valid,
      outs_ready(0) => fork7_outs_0_ready,
      outs_ready(1) => fork7_outs_1_ready,
      outs_ready(2) => fork7_outs_2_ready
    );

  buffer119 : entity work.handshake_buffer_1(arch)
    port map(
      ins => fork6_outs_1,
      ins_valid => fork6_outs_1_valid,
      ins_ready => fork6_outs_1_ready,
      clk => clk,
      rst => rst,
      outs => buffer119_outs,
      outs_valid => buffer119_outs_valid,
      outs_ready => buffer119_outs_ready
    );

  buffer120 : entity work.handshake_buffer_1(arch)
    port map(
      ins => buffer119_outs,
      ins_valid => buffer119_outs_valid,
      ins_ready => buffer119_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer120_outs,
      outs_valid => buffer120_outs_valid,
      outs_ready => buffer120_outs_ready
    );

  buffer121 : entity work.handshake_buffer_1(arch)
    port map(
      ins => buffer120_outs,
      ins_valid => buffer120_outs_valid,
      ins_ready => buffer120_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer121_outs,
      outs_valid => buffer121_outs_valid,
      outs_ready => buffer121_outs_ready
    );

  buffer122 : entity work.handshake_buffer_1(arch)
    port map(
      ins => buffer121_outs,
      ins_valid => buffer121_outs_valid,
      ins_ready => buffer121_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer122_outs,
      outs_valid => buffer122_outs_valid,
      outs_ready => buffer122_outs_ready
    );

  buffer123 : entity work.handshake_buffer_1(arch)
    port map(
      ins => buffer122_outs,
      ins_valid => buffer122_outs_valid,
      ins_ready => buffer122_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer123_outs,
      outs_valid => buffer123_outs_valid,
      outs_ready => buffer123_outs_ready
    );

  mux8 : entity work.handshake_mux_2(arch)
    port map(
      index => buffer123_outs,
      index_valid => buffer123_outs_valid,
      index_ready => buffer123_outs_ready,
      ins(0) => extsi9_outs,
      ins(1) => cond_br17_trueOut,
      ins_valid(0) => extsi9_outs_valid,
      ins_valid(1) => cond_br17_trueOut_valid,
      ins_ready(0) => extsi9_outs_ready,
      ins_ready(1) => cond_br17_trueOut_ready,
      clk => clk,
      rst => rst,
      outs => mux8_outs,
      outs_valid => mux8_outs_valid,
      outs_ready => mux8_outs_ready
    );

  buffer114 : entity work.handshake_buffer_1(arch)
    port map(
      ins => fork6_outs_0,
      ins_valid => fork6_outs_0_valid,
      ins_ready => fork6_outs_0_ready,
      clk => clk,
      rst => rst,
      outs => buffer114_outs,
      outs_valid => buffer114_outs_valid,
      outs_ready => buffer114_outs_ready
    );

  buffer115 : entity work.handshake_buffer_1(arch)
    port map(
      ins => buffer114_outs,
      ins_valid => buffer114_outs_valid,
      ins_ready => buffer114_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer115_outs,
      outs_valid => buffer115_outs_valid,
      outs_ready => buffer115_outs_ready
    );

  buffer116 : entity work.handshake_buffer_1(arch)
    port map(
      ins => buffer115_outs,
      ins_valid => buffer115_outs_valid,
      ins_ready => buffer115_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer116_outs,
      outs_valid => buffer116_outs_valid,
      outs_ready => buffer116_outs_ready
    );

  buffer117 : entity work.handshake_buffer_1(arch)
    port map(
      ins => buffer116_outs,
      ins_valid => buffer116_outs_valid,
      ins_ready => buffer116_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer117_outs,
      outs_valid => buffer117_outs_valid,
      outs_ready => buffer117_outs_ready
    );

  buffer118 : entity work.handshake_buffer_1(arch)
    port map(
      ins => buffer117_outs,
      ins_valid => buffer117_outs_valid,
      ins_ready => buffer117_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer118_outs,
      outs_valid => buffer118_outs_valid,
      outs_ready => buffer118_outs_ready
    );

  mux9 : entity work.handshake_mux_1(arch)
    port map(
      index => buffer118_outs,
      index_valid => buffer118_outs_valid,
      index_ready => buffer118_outs_ready,
      ins(0) => extsi10_outs,
      ins(1) => cond_br18_trueOut,
      ins_valid(0) => extsi10_outs_valid,
      ins_valid(1) => cond_br18_trueOut_valid,
      ins_ready(0) => extsi10_outs_ready,
      ins_ready(1) => cond_br18_trueOut_ready,
      clk => clk,
      rst => rst,
      outs => mux9_outs,
      outs_valid => mux9_outs_valid,
      outs_ready => mux9_outs_ready
    );

  buffer145 : entity work.handshake_buffer_3(arch)
    port map(
      ins => mux9_outs,
      ins_valid => mux9_outs_valid,
      ins_ready => mux9_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer145_outs,
      outs_valid => buffer145_outs_valid,
      outs_ready => buffer145_outs_ready
    );

  buffer146 : entity work.handshake_buffer_4(arch)
    port map(
      ins => buffer145_outs,
      ins_valid => buffer145_outs_valid,
      ins_ready => buffer145_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer146_outs,
      outs_valid => buffer146_outs_valid,
      outs_ready => buffer146_outs_ready
    );

  buffer147 : entity work.handshake_buffer_4(arch)
    port map(
      ins => buffer146_outs,
      ins_valid => buffer146_outs_valid,
      ins_ready => buffer146_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer147_outs,
      outs_valid => buffer147_outs_valid,
      outs_ready => buffer147_outs_ready
    );

  buffer148 : entity work.handshake_buffer_4(arch)
    port map(
      ins => buffer147_outs,
      ins_valid => buffer147_outs_valid,
      ins_ready => buffer147_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer148_outs,
      outs_valid => buffer148_outs_valid,
      outs_ready => buffer148_outs_ready
    );

  buffer149 : entity work.handshake_buffer_4(arch)
    port map(
      ins => buffer148_outs,
      ins_valid => buffer148_outs_valid,
      ins_ready => buffer148_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer149_outs,
      outs_valid => buffer149_outs_valid,
      outs_ready => buffer149_outs_ready
    );

  buffer150 : entity work.handshake_buffer_4(arch)
    port map(
      ins => buffer149_outs,
      ins_valid => buffer149_outs_valid,
      ins_ready => buffer149_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer150_outs,
      outs_valid => buffer150_outs_valid,
      outs_ready => buffer150_outs_ready
    );

  fork8 : entity work.handshake_fork_5(arch)
    port map(
      ins => buffer150_outs,
      ins_valid => buffer150_outs_valid,
      ins_ready => buffer150_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork8_outs_0,
      outs(1) => fork8_outs_1,
      outs_valid(0) => fork8_outs_0_valid,
      outs_valid(1) => fork8_outs_1_valid,
      outs_ready(0) => fork8_outs_0_ready,
      outs_ready(1) => fork8_outs_1_ready
    );

  buffer156 : entity work.handshake_buffer_4(arch)
    port map(
      ins => fork8_outs_1,
      ins_valid => fork8_outs_1_valid,
      ins_ready => fork8_outs_1_ready,
      clk => clk,
      rst => rst,
      outs => buffer156_outs,
      outs_valid => buffer156_outs_valid,
      outs_ready => buffer156_outs_ready
    );

  buffer157 : entity work.handshake_buffer_4(arch)
    port map(
      ins => buffer156_outs,
      ins_valid => buffer156_outs_valid,
      ins_ready => buffer156_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer157_outs,
      outs_valid => buffer157_outs_valid,
      outs_ready => buffer157_outs_ready
    );

  buffer158 : entity work.handshake_buffer_4(arch)
    port map(
      ins => buffer157_outs,
      ins_valid => buffer157_outs_valid,
      ins_ready => buffer157_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer158_outs,
      outs_valid => buffer158_outs_valid,
      outs_ready => buffer158_outs_ready
    );

  buffer159 : entity work.handshake_buffer_4(arch)
    port map(
      ins => buffer158_outs,
      ins_valid => buffer158_outs_valid,
      ins_ready => buffer158_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer159_outs,
      outs_valid => buffer159_outs_valid,
      outs_ready => buffer159_outs_ready
    );

  buffer160 : entity work.handshake_buffer_4(arch)
    port map(
      ins => buffer159_outs,
      ins_valid => buffer159_outs_valid,
      ins_ready => buffer159_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer160_outs,
      outs_valid => buffer160_outs_valid,
      outs_ready => buffer160_outs_ready
    );

  extsi11 : entity work.handshake_extsi_1(arch)
    port map(
      ins => buffer160_outs,
      ins_valid => buffer160_outs_valid,
      ins_ready => buffer160_outs_ready,
      clk => clk,
      rst => rst,
      outs => extsi11_outs,
      outs_valid => extsi11_outs_valid,
      outs_ready => extsi11_outs_ready
    );

  buffer151 : entity work.handshake_buffer_4(arch)
    port map(
      ins => fork8_outs_0,
      ins_valid => fork8_outs_0_valid,
      ins_ready => fork8_outs_0_ready,
      clk => clk,
      rst => rst,
      outs => buffer151_outs,
      outs_valid => buffer151_outs_valid,
      outs_ready => buffer151_outs_ready
    );

  buffer152 : entity work.handshake_buffer_4(arch)
    port map(
      ins => buffer151_outs,
      ins_valid => buffer151_outs_valid,
      ins_ready => buffer151_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer152_outs,
      outs_valid => buffer152_outs_valid,
      outs_ready => buffer152_outs_ready
    );

  buffer153 : entity work.handshake_buffer_4(arch)
    port map(
      ins => buffer152_outs,
      ins_valid => buffer152_outs_valid,
      ins_ready => buffer152_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer153_outs,
      outs_valid => buffer153_outs_valid,
      outs_ready => buffer153_outs_ready
    );

  buffer154 : entity work.handshake_buffer_4(arch)
    port map(
      ins => buffer153_outs,
      ins_valid => buffer153_outs_valid,
      ins_ready => buffer153_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer154_outs,
      outs_valid => buffer154_outs_valid,
      outs_ready => buffer154_outs_ready
    );

  buffer155 : entity work.handshake_buffer_4(arch)
    port map(
      ins => buffer154_outs,
      ins_valid => buffer154_outs_valid,
      ins_ready => buffer154_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer155_outs,
      outs_valid => buffer155_outs_valid,
      outs_ready => buffer155_outs_ready
    );

  extsi12 : entity work.handshake_extsi_2(arch)
    port map(
      ins => buffer155_outs,
      ins_valid => buffer155_outs_valid,
      ins_ready => buffer155_outs_ready,
      clk => clk,
      rst => rst,
      outs => extsi12_outs,
      outs_valid => extsi12_outs_valid,
      outs_ready => extsi12_outs_ready
    );

  buffer129 : entity work.handshake_buffer_0(arch)
    port map(
      ins_valid => fork7_outs_1_valid,
      ins_ready => fork7_outs_1_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer129_outs_valid,
      outs_ready => buffer129_outs_ready
    );

  buffer130 : entity work.handshake_buffer_0(arch)
    port map(
      ins_valid => buffer129_outs_valid,
      ins_ready => buffer129_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer130_outs_valid,
      outs_ready => buffer130_outs_ready
    );

  buffer131 : entity work.handshake_buffer_0(arch)
    port map(
      ins_valid => buffer130_outs_valid,
      ins_ready => buffer130_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer131_outs_valid,
      outs_ready => buffer131_outs_ready
    );

  buffer132 : entity work.handshake_buffer_0(arch)
    port map(
      ins_valid => buffer131_outs_valid,
      ins_ready => buffer131_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer132_outs_valid,
      outs_ready => buffer132_outs_ready
    );

  buffer133 : entity work.handshake_buffer_0(arch)
    port map(
      ins_valid => buffer132_outs_valid,
      ins_ready => buffer132_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer133_outs_valid,
      outs_ready => buffer133_outs_ready
    );

  constant9 : entity work.handshake_constant_1(arch)
    port map(
      ctrl_valid => buffer133_outs_valid,
      ctrl_ready => buffer133_outs_ready,
      clk => clk,
      rst => rst,
      outs => constant9_outs,
      outs_valid => constant9_outs_valid,
      outs_ready => constant9_outs_ready
    );

  extsi13 : entity work.handshake_extsi_1(arch)
    port map(
      ins => constant9_outs,
      ins_valid => constant9_outs_valid,
      ins_ready => constant9_outs_ready,
      clk => clk,
      rst => rst,
      outs => extsi13_outs,
      outs_valid => extsi13_outs_valid,
      outs_ready => extsi13_outs_ready
    );

  buffer124 : entity work.handshake_buffer_0(arch)
    port map(
      ins_valid => fork7_outs_0_valid,
      ins_ready => fork7_outs_0_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer124_outs_valid,
      outs_ready => buffer124_outs_ready
    );

  buffer125 : entity work.handshake_buffer_0(arch)
    port map(
      ins_valid => buffer124_outs_valid,
      ins_ready => buffer124_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer125_outs_valid,
      outs_ready => buffer125_outs_ready
    );

  buffer126 : entity work.handshake_buffer_0(arch)
    port map(
      ins_valid => buffer125_outs_valid,
      ins_ready => buffer125_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer126_outs_valid,
      outs_ready => buffer126_outs_ready
    );

  buffer127 : entity work.handshake_buffer_0(arch)
    port map(
      ins_valid => buffer126_outs_valid,
      ins_ready => buffer126_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer127_outs_valid,
      outs_ready => buffer127_outs_ready
    );

  buffer128 : entity work.handshake_buffer_0(arch)
    port map(
      ins_valid => buffer127_outs_valid,
      ins_ready => buffer127_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer128_outs_valid,
      outs_ready => buffer128_outs_ready
    );

  constant10 : entity work.handshake_constant_2(arch)
    port map(
      ctrl_valid => buffer128_outs_valid,
      ctrl_ready => buffer128_outs_ready,
      clk => clk,
      rst => rst,
      outs => constant10_outs,
      outs_valid => constant10_outs_valid,
      outs_ready => constant10_outs_ready
    );

  extsi14 : entity work.handshake_extsi_3(arch)
    port map(
      ins => constant10_outs,
      ins_valid => constant10_outs_valid,
      ins_ready => constant10_outs_ready,
      clk => clk,
      rst => rst,
      outs => extsi14_outs,
      outs_valid => extsi14_outs_valid,
      outs_ready => extsi14_outs_ready
    );

  buffer139 : entity work.handshake_buffer_5(arch)
    port map(
      ins => mux8_outs,
      ins_valid => mux8_outs_valid,
      ins_ready => mux8_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer139_outs,
      outs_valid => buffer139_outs_valid,
      outs_ready => buffer139_outs_ready
    );

  buffer140 : entity work.handshake_buffer_6(arch)
    port map(
      ins => buffer139_outs,
      ins_valid => buffer139_outs_valid,
      ins_ready => buffer139_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer140_outs,
      outs_valid => buffer140_outs_valid,
      outs_ready => buffer140_outs_ready
    );

  buffer141 : entity work.handshake_buffer_6(arch)
    port map(
      ins => buffer140_outs,
      ins_valid => buffer140_outs_valid,
      ins_ready => buffer140_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer141_outs,
      outs_valid => buffer141_outs_valid,
      outs_ready => buffer141_outs_ready
    );

  buffer142 : entity work.handshake_buffer_6(arch)
    port map(
      ins => buffer141_outs,
      ins_valid => buffer141_outs_valid,
      ins_ready => buffer141_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer142_outs,
      outs_valid => buffer142_outs_valid,
      outs_ready => buffer142_outs_ready
    );

  buffer143 : entity work.handshake_buffer_6(arch)
    port map(
      ins => buffer142_outs,
      ins_valid => buffer142_outs_valid,
      ins_ready => buffer142_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer143_outs,
      outs_valid => buffer143_outs_valid,
      outs_ready => buffer143_outs_ready
    );

  buffer144 : entity work.handshake_buffer_6(arch)
    port map(
      ins => buffer143_outs,
      ins_valid => buffer143_outs_valid,
      ins_ready => buffer143_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer144_outs,
      outs_valid => buffer144_outs_valid,
      outs_ready => buffer144_outs_ready
    );

  muli0 : entity work.handshake_muli_0(arch)
    port map(
      lhs => buffer144_outs,
      lhs_valid => buffer144_outs_valid,
      lhs_ready => buffer144_outs_ready,
      rhs => extsi12_outs,
      rhs_valid => extsi12_outs_valid,
      rhs_ready => extsi12_outs_ready,
      clk => clk,
      rst => rst,
      result => muli0_result,
      result_valid => muli0_result_valid,
      result_ready => muli0_result_ready
    );

  addi1 : entity work.handshake_addi_0(arch)
    port map(
      lhs => extsi11_outs,
      lhs_valid => extsi11_outs_valid,
      lhs_ready => extsi11_outs_ready,
      rhs => extsi14_outs,
      rhs_valid => extsi14_outs_valid,
      rhs_ready => extsi14_outs_ready,
      clk => clk,
      rst => rst,
      result => addi1_result,
      result_valid => addi1_result_valid,
      result_ready => addi1_result_ready
    );

  fork9 : entity work.handshake_fork_6(arch)
    port map(
      ins => addi1_result,
      ins_valid => addi1_result_valid,
      ins_ready => addi1_result_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork9_outs_0,
      outs(1) => fork9_outs_1,
      outs_valid(0) => fork9_outs_0_valid,
      outs_valid(1) => fork9_outs_1_valid,
      outs_ready(0) => fork9_outs_0_ready,
      outs_ready(1) => fork9_outs_1_ready
    );

  buffer166 : entity work.handshake_buffer_7(arch)
    port map(
      ins => fork9_outs_1,
      ins_valid => fork9_outs_1_valid,
      ins_ready => fork9_outs_1_ready,
      clk => clk,
      rst => rst,
      outs => buffer166_outs,
      outs_valid => buffer166_outs_valid,
      outs_ready => buffer166_outs_ready
    );

  buffer167 : entity work.handshake_buffer_7(arch)
    port map(
      ins => buffer166_outs,
      ins_valid => buffer166_outs_valid,
      ins_ready => buffer166_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer167_outs,
      outs_valid => buffer167_outs_valid,
      outs_ready => buffer167_outs_ready
    );

  buffer168 : entity work.handshake_buffer_7(arch)
    port map(
      ins => buffer167_outs,
      ins_valid => buffer167_outs_valid,
      ins_ready => buffer167_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer168_outs,
      outs_valid => buffer168_outs_valid,
      outs_ready => buffer168_outs_ready
    );

  buffer169 : entity work.handshake_buffer_7(arch)
    port map(
      ins => buffer168_outs,
      ins_valid => buffer168_outs_valid,
      ins_ready => buffer168_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer169_outs,
      outs_valid => buffer169_outs_valid,
      outs_ready => buffer169_outs_ready
    );

  buffer170 : entity work.handshake_buffer_7(arch)
    port map(
      ins => buffer169_outs,
      ins_valid => buffer169_outs_valid,
      ins_ready => buffer169_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer170_outs,
      outs_valid => buffer170_outs_valid,
      outs_ready => buffer170_outs_ready
    );

  trunci1 : entity work.handshake_trunci_1(arch)
    port map(
      ins => buffer170_outs,
      ins_valid => buffer170_outs_valid,
      ins_ready => buffer170_outs_ready,
      clk => clk,
      rst => rst,
      outs => trunci1_outs,
      outs_valid => trunci1_outs_valid,
      outs_ready => trunci1_outs_ready
    );

  buffer161 : entity work.handshake_buffer_7(arch)
    port map(
      ins => fork9_outs_0,
      ins_valid => fork9_outs_0_valid,
      ins_ready => fork9_outs_0_ready,
      clk => clk,
      rst => rst,
      outs => buffer161_outs,
      outs_valid => buffer161_outs_valid,
      outs_ready => buffer161_outs_ready
    );

  buffer162 : entity work.handshake_buffer_7(arch)
    port map(
      ins => buffer161_outs,
      ins_valid => buffer161_outs_valid,
      ins_ready => buffer161_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer162_outs,
      outs_valid => buffer162_outs_valid,
      outs_ready => buffer162_outs_ready
    );

  buffer163 : entity work.handshake_buffer_7(arch)
    port map(
      ins => buffer162_outs,
      ins_valid => buffer162_outs_valid,
      ins_ready => buffer162_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer163_outs,
      outs_valid => buffer163_outs_valid,
      outs_ready => buffer163_outs_ready
    );

  buffer164 : entity work.handshake_buffer_7(arch)
    port map(
      ins => buffer163_outs,
      ins_valid => buffer163_outs_valid,
      ins_ready => buffer163_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer164_outs,
      outs_valid => buffer164_outs_valid,
      outs_ready => buffer164_outs_ready
    );

  buffer165 : entity work.handshake_buffer_7(arch)
    port map(
      ins => buffer164_outs,
      ins_valid => buffer164_outs_valid,
      ins_ready => buffer164_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer165_outs,
      outs_valid => buffer165_outs_valid,
      outs_ready => buffer165_outs_ready
    );

  cmpi0 : entity work.handshake_cmpi_0(arch)
    port map(
      lhs => buffer165_outs,
      lhs_valid => buffer165_outs_valid,
      lhs_ready => buffer165_outs_ready,
      rhs => extsi13_outs,
      rhs_valid => extsi13_outs_valid,
      rhs_ready => extsi13_outs_ready,
      clk => clk,
      rst => rst,
      result => cmpi0_result,
      result_valid => cmpi0_result_valid,
      result_ready => cmpi0_result_ready
    );

  fork10 : entity work.handshake_fork_7(arch)
    port map(
      ins => cmpi0_result,
      ins_valid => cmpi0_result_valid,
      ins_ready => cmpi0_result_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork10_outs_0,
      outs(1) => fork10_outs_1,
      outs(2) => fork10_outs_2,
      outs_valid(0) => fork10_outs_0_valid,
      outs_valid(1) => fork10_outs_1_valid,
      outs_valid(2) => fork10_outs_2_valid,
      outs_ready(0) => fork10_outs_0_ready,
      outs_ready(1) => fork10_outs_1_ready,
      outs_ready(2) => fork10_outs_2_ready
    );

  buffer103 : entity work.handshake_buffer_6(arch)
    port map(
      ins => fork5_outs_1,
      ins_valid => fork5_outs_1_valid,
      ins_ready => fork5_outs_1_ready,
      clk => clk,
      rst => rst,
      outs => buffer103_outs,
      outs_valid => buffer103_outs_valid,
      outs_ready => buffer103_outs_ready
    );

  buffer104 : entity work.handshake_buffer_6(arch)
    port map(
      ins => buffer103_outs,
      ins_valid => buffer103_outs_valid,
      ins_ready => buffer103_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer104_outs,
      outs_valid => buffer104_outs_valid,
      outs_ready => buffer104_outs_ready
    );

  buffer105 : entity work.handshake_buffer_6(arch)
    port map(
      ins => buffer104_outs,
      ins_valid => buffer104_outs_valid,
      ins_ready => buffer104_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer105_outs,
      outs_valid => buffer105_outs_valid,
      outs_ready => buffer105_outs_ready
    );

  buffer106 : entity work.handshake_buffer_6(arch)
    port map(
      ins => buffer105_outs,
      ins_valid => buffer105_outs_valid,
      ins_ready => buffer105_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer106_outs,
      outs_valid => buffer106_outs_valid,
      outs_ready => buffer106_outs_ready
    );

  buffer107 : entity work.handshake_buffer_6(arch)
    port map(
      ins => buffer106_outs,
      ins_valid => buffer106_outs_valid,
      ins_ready => buffer106_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer107_outs,
      outs_valid => buffer107_outs_valid,
      outs_ready => buffer107_outs_ready
    );

  buffer201 : entity work.handshake_buffer_1(arch)
    port map(
      ins => fork12_outs_1,
      ins_valid => fork12_outs_1_valid,
      ins_ready => fork12_outs_1_ready,
      clk => clk,
      rst => rst,
      outs => buffer201_outs,
      outs_valid => buffer201_outs_valid,
      outs_ready => buffer201_outs_ready
    );

  buffer202 : entity work.handshake_buffer_1(arch)
    port map(
      ins => buffer201_outs,
      ins_valid => buffer201_outs_valid,
      ins_ready => buffer201_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer202_outs,
      outs_valid => buffer202_outs_valid,
      outs_ready => buffer202_outs_ready
    );

  buffer203 : entity work.handshake_buffer_1(arch)
    port map(
      ins => buffer202_outs,
      ins_valid => buffer202_outs_valid,
      ins_ready => buffer202_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer203_outs,
      outs_valid => buffer203_outs_valid,
      outs_ready => buffer203_outs_ready
    );

  buffer204 : entity work.handshake_buffer_1(arch)
    port map(
      ins => buffer203_outs,
      ins_valid => buffer203_outs_valid,
      ins_ready => buffer203_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer204_outs,
      outs_valid => buffer204_outs_valid,
      outs_ready => buffer204_outs_ready
    );

  buffer205 : entity work.handshake_buffer_1(arch)
    port map(
      ins => buffer204_outs,
      ins_valid => buffer204_outs_valid,
      ins_ready => buffer204_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer205_outs,
      outs_valid => buffer205_outs_valid,
      outs_ready => buffer205_outs_ready
    );

  cond_br20 : entity work.handshake_cond_br_0(arch)
    port map(
      condition => buffer205_outs,
      condition_valid => buffer205_outs_valid,
      condition_ready => buffer205_outs_ready,
      data => buffer107_outs,
      data_valid => buffer107_outs_valid,
      data_ready => buffer107_outs_ready,
      clk => clk,
      rst => rst,
      trueOut => cond_br20_trueOut,
      trueOut_valid => cond_br20_trueOut_valid,
      trueOut_ready => cond_br20_trueOut_ready,
      falseOut => cond_br20_falseOut,
      falseOut_valid => cond_br20_falseOut_valid,
      falseOut_ready => cond_br20_falseOut_ready
    );

  sink2 : entity work.handshake_sink_2(arch)
    port map(
      ins => cond_br20_trueOut,
      ins_valid => cond_br20_trueOut_valid,
      ins_ready => cond_br20_trueOut_ready,
      clk => clk,
      rst => rst
    );

  buffer206 : entity work.handshake_buffer_1(arch)
    port map(
      ins => fork12_outs_2,
      ins_valid => fork12_outs_2_valid,
      ins_ready => fork12_outs_2_ready,
      clk => clk,
      rst => rst,
      outs => buffer206_outs,
      outs_valid => buffer206_outs_valid,
      outs_ready => buffer206_outs_ready
    );

  buffer207 : entity work.handshake_buffer_1(arch)
    port map(
      ins => buffer206_outs,
      ins_valid => buffer206_outs_valid,
      ins_ready => buffer206_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer207_outs,
      outs_valid => buffer207_outs_valid,
      outs_ready => buffer207_outs_ready
    );

  buffer208 : entity work.handshake_buffer_1(arch)
    port map(
      ins => buffer207_outs,
      ins_valid => buffer207_outs_valid,
      ins_ready => buffer207_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer208_outs,
      outs_valid => buffer208_outs_valid,
      outs_ready => buffer208_outs_ready
    );

  buffer209 : entity work.handshake_buffer_1(arch)
    port map(
      ins => buffer208_outs,
      ins_valid => buffer208_outs_valid,
      ins_ready => buffer208_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer209_outs,
      outs_valid => buffer209_outs_valid,
      outs_ready => buffer209_outs_ready
    );

  buffer210 : entity work.handshake_buffer_1(arch)
    port map(
      ins => buffer209_outs,
      ins_valid => buffer209_outs_valid,
      ins_ready => buffer209_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer210_outs,
      outs_valid => buffer210_outs_valid,
      outs_ready => buffer210_outs_ready
    );

  cond_br21 : entity work.handshake_cond_br_1(arch)
    port map(
      condition => buffer210_outs,
      condition_valid => buffer210_outs_valid,
      condition_ready => buffer210_outs_ready,
      data => trunci2_outs,
      data_valid => trunci2_outs_valid,
      data_ready => trunci2_outs_ready,
      clk => clk,
      rst => rst,
      trueOut => cond_br21_trueOut,
      trueOut_valid => cond_br21_trueOut_valid,
      trueOut_ready => cond_br21_trueOut_ready,
      falseOut => cond_br21_falseOut,
      falseOut_valid => cond_br21_falseOut_valid,
      falseOut_ready => cond_br21_falseOut_ready
    );

  sink3 : entity work.handshake_sink_0(arch)
    port map(
      ins => cond_br21_falseOut,
      ins_valid => cond_br21_falseOut_valid,
      ins_ready => cond_br21_falseOut_ready,
      clk => clk,
      rst => rst
    );

  buffer62 : entity work.handshake_buffer_0(arch)
    port map(
      ins_valid => fork3_outs_2_valid,
      ins_ready => fork3_outs_2_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer62_outs_valid,
      outs_ready => buffer62_outs_ready
    );

  buffer63 : entity work.handshake_buffer_0(arch)
    port map(
      ins_valid => buffer62_outs_valid,
      ins_ready => buffer62_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer63_outs_valid,
      outs_ready => buffer63_outs_ready
    );

  buffer64 : entity work.handshake_buffer_0(arch)
    port map(
      ins_valid => buffer63_outs_valid,
      ins_ready => buffer63_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer64_outs_valid,
      outs_ready => buffer64_outs_ready
    );

  buffer65 : entity work.handshake_buffer_0(arch)
    port map(
      ins_valid => buffer64_outs_valid,
      ins_ready => buffer64_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer65_outs_valid,
      outs_ready => buffer65_outs_ready
    );

  buffer66 : entity work.handshake_buffer_0(arch)
    port map(
      ins_valid => buffer65_outs_valid,
      ins_ready => buffer65_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer66_outs_valid,
      outs_ready => buffer66_outs_ready
    );

  buffer211 : entity work.handshake_buffer_1(arch)
    port map(
      ins => fork12_outs_3,
      ins_valid => fork12_outs_3_valid,
      ins_ready => fork12_outs_3_ready,
      clk => clk,
      rst => rst,
      outs => buffer211_outs,
      outs_valid => buffer211_outs_valid,
      outs_ready => buffer211_outs_ready
    );

  buffer212 : entity work.handshake_buffer_1(arch)
    port map(
      ins => buffer211_outs,
      ins_valid => buffer211_outs_valid,
      ins_ready => buffer211_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer212_outs,
      outs_valid => buffer212_outs_valid,
      outs_ready => buffer212_outs_ready
    );

  buffer213 : entity work.handshake_buffer_1(arch)
    port map(
      ins => buffer212_outs,
      ins_valid => buffer212_outs_valid,
      ins_ready => buffer212_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer213_outs,
      outs_valid => buffer213_outs_valid,
      outs_ready => buffer213_outs_ready
    );

  buffer214 : entity work.handshake_buffer_1(arch)
    port map(
      ins => buffer213_outs,
      ins_valid => buffer213_outs_valid,
      ins_ready => buffer213_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer214_outs,
      outs_valid => buffer214_outs_valid,
      outs_ready => buffer214_outs_ready
    );

  buffer215 : entity work.handshake_buffer_1(arch)
    port map(
      ins => buffer214_outs,
      ins_valid => buffer214_outs_valid,
      ins_ready => buffer214_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer215_outs,
      outs_valid => buffer215_outs_valid,
      outs_ready => buffer215_outs_ready
    );

  cond_br22 : entity work.handshake_cond_br_2(arch)
    port map(
      condition => buffer215_outs,
      condition_valid => buffer215_outs_valid,
      condition_ready => buffer215_outs_ready,
      data_valid => buffer66_outs_valid,
      data_ready => buffer66_outs_ready,
      clk => clk,
      rst => rst,
      trueOut_valid => cond_br22_trueOut_valid,
      trueOut_ready => cond_br22_trueOut_ready,
      falseOut_valid => cond_br22_falseOut_valid,
      falseOut_ready => cond_br22_falseOut_ready
    );

  sink4 : entity work.handshake_sink_1(arch)
    port map(
      ins_valid => cond_br22_falseOut_valid,
      ins_ready => cond_br22_falseOut_ready,
      clk => clk,
      rst => rst
    );

  buffer5 : entity work.handshake_buffer_0(arch)
    port map(
      ins_valid => fork0_outs_1_valid,
      ins_ready => fork0_outs_1_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer5_outs_valid,
      outs_ready => buffer5_outs_ready
    );

  buffer6 : entity work.handshake_buffer_0(arch)
    port map(
      ins_valid => buffer5_outs_valid,
      ins_ready => buffer5_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer6_outs_valid,
      outs_ready => buffer6_outs_ready
    );

  buffer7 : entity work.handshake_buffer_0(arch)
    port map(
      ins_valid => buffer6_outs_valid,
      ins_ready => buffer6_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer7_outs_valid,
      outs_ready => buffer7_outs_ready
    );

  buffer8 : entity work.handshake_buffer_0(arch)
    port map(
      ins_valid => buffer7_outs_valid,
      ins_ready => buffer7_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer8_outs_valid,
      outs_ready => buffer8_outs_ready
    );

  buffer9 : entity work.handshake_buffer_0(arch)
    port map(
      ins_valid => buffer8_outs_valid,
      ins_ready => buffer8_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer9_outs_valid,
      outs_ready => buffer9_outs_ready
    );

  constant11 : entity work.handshake_constant_2(arch)
    port map(
      ctrl_valid => buffer9_outs_valid,
      ctrl_ready => buffer9_outs_ready,
      clk => clk,
      rst => rst,
      outs => constant11_outs,
      outs_valid => constant11_outs_valid,
      outs_ready => constant11_outs_ready
    );

  extsi4 : entity work.handshake_extsi_4(arch)
    port map(
      ins => constant11_outs,
      ins_valid => constant11_outs_valid,
      ins_ready => constant11_outs_ready,
      clk => clk,
      rst => rst,
      outs => extsi4_outs,
      outs_valid => extsi4_outs_valid,
      outs_ready => extsi4_outs_ready
    );

  buffer57 : entity work.handshake_buffer_0(arch)
    port map(
      ins_valid => fork3_outs_1_valid,
      ins_ready => fork3_outs_1_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer57_outs_valid,
      outs_ready => buffer57_outs_ready
    );

  buffer58 : entity work.handshake_buffer_0(arch)
    port map(
      ins_valid => buffer57_outs_valid,
      ins_ready => buffer57_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer58_outs_valid,
      outs_ready => buffer58_outs_ready
    );

  buffer59 : entity work.handshake_buffer_0(arch)
    port map(
      ins_valid => buffer58_outs_valid,
      ins_ready => buffer58_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer59_outs_valid,
      outs_ready => buffer59_outs_ready
    );

  buffer60 : entity work.handshake_buffer_0(arch)
    port map(
      ins_valid => buffer59_outs_valid,
      ins_ready => buffer59_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer60_outs_valid,
      outs_ready => buffer60_outs_ready
    );

  buffer61 : entity work.handshake_buffer_0(arch)
    port map(
      ins_valid => buffer60_outs_valid,
      ins_ready => buffer60_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer61_outs_valid,
      outs_ready => buffer61_outs_ready
    );

  constant13 : entity work.handshake_constant_1(arch)
    port map(
      ctrl_valid => buffer61_outs_valid,
      ctrl_ready => buffer61_outs_ready,
      clk => clk,
      rst => rst,
      outs => constant13_outs,
      outs_valid => constant13_outs_valid,
      outs_ready => constant13_outs_ready
    );

  extsi15 : entity work.handshake_extsi_1(arch)
    port map(
      ins => constant13_outs,
      ins_valid => constant13_outs_valid,
      ins_ready => constant13_outs_ready,
      clk => clk,
      rst => rst,
      outs => extsi15_outs,
      outs_valid => extsi15_outs_valid,
      outs_ready => extsi15_outs_ready
    );

  buffer52 : entity work.handshake_buffer_0(arch)
    port map(
      ins_valid => fork3_outs_0_valid,
      ins_ready => fork3_outs_0_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer52_outs_valid,
      outs_ready => buffer52_outs_ready
    );

  buffer53 : entity work.handshake_buffer_0(arch)
    port map(
      ins_valid => buffer52_outs_valid,
      ins_ready => buffer52_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer53_outs_valid,
      outs_ready => buffer53_outs_ready
    );

  buffer54 : entity work.handshake_buffer_0(arch)
    port map(
      ins_valid => buffer53_outs_valid,
      ins_ready => buffer53_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer54_outs_valid,
      outs_ready => buffer54_outs_ready
    );

  buffer55 : entity work.handshake_buffer_0(arch)
    port map(
      ins_valid => buffer54_outs_valid,
      ins_ready => buffer54_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer55_outs_valid,
      outs_ready => buffer55_outs_ready
    );

  buffer56 : entity work.handshake_buffer_0(arch)
    port map(
      ins_valid => buffer55_outs_valid,
      ins_ready => buffer55_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer56_outs_valid,
      outs_ready => buffer56_outs_ready
    );

  constant14 : entity work.handshake_constant_2(arch)
    port map(
      ctrl_valid => buffer56_outs_valid,
      ctrl_ready => buffer56_outs_ready,
      clk => clk,
      rst => rst,
      outs => constant14_outs,
      outs_valid => constant14_outs_valid,
      outs_ready => constant14_outs_ready
    );

  extsi16 : entity work.handshake_extsi_3(arch)
    port map(
      ins => constant14_outs,
      ins_valid => constant14_outs_valid,
      ins_ready => constant14_outs_ready,
      clk => clk,
      rst => rst,
      outs => extsi16_outs,
      outs_valid => extsi16_outs_valid,
      outs_ready => extsi16_outs_ready
    );

  buffer98 : entity work.handshake_buffer_6(arch)
    port map(
      ins => fork5_outs_0,
      ins_valid => fork5_outs_0_valid,
      ins_ready => fork5_outs_0_ready,
      clk => clk,
      rst => rst,
      outs => buffer98_outs,
      outs_valid => buffer98_outs_valid,
      outs_ready => buffer98_outs_ready
    );

  buffer99 : entity work.handshake_buffer_6(arch)
    port map(
      ins => buffer98_outs,
      ins_valid => buffer98_outs_valid,
      ins_ready => buffer98_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer99_outs,
      outs_valid => buffer99_outs_valid,
      outs_ready => buffer99_outs_ready
    );

  buffer100 : entity work.handshake_buffer_6(arch)
    port map(
      ins => buffer99_outs,
      ins_valid => buffer99_outs_valid,
      ins_ready => buffer99_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer100_outs,
      outs_valid => buffer100_outs_valid,
      outs_ready => buffer100_outs_ready
    );

  buffer101 : entity work.handshake_buffer_6(arch)
    port map(
      ins => buffer100_outs,
      ins_valid => buffer100_outs_valid,
      ins_ready => buffer100_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer101_outs,
      outs_valid => buffer101_outs_valid,
      outs_ready => buffer101_outs_ready
    );

  buffer102 : entity work.handshake_buffer_6(arch)
    port map(
      ins => buffer101_outs,
      ins_valid => buffer101_outs_valid,
      ins_ready => buffer101_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer102_outs,
      outs_valid => buffer102_outs_valid,
      outs_ready => buffer102_outs_ready
    );

  store0 : entity work.handshake_store_0(arch)
    port map(
      addrIn => trunci0_outs,
      addrIn_valid => trunci0_outs_valid,
      addrIn_ready => trunci0_outs_ready,
      dataIn => buffer102_outs,
      dataIn_valid => buffer102_outs_valid,
      dataIn_ready => buffer102_outs_ready,
      clk => clk,
      rst => rst,
      addrOut => store0_addrOut,
      addrOut_valid => store0_addrOut_valid,
      addrOut_ready => store0_addrOut_ready,
      dataToMem => store0_dataToMem,
      dataToMem_valid => store0_dataToMem_valid,
      dataToMem_ready => store0_dataToMem_ready
    );

  addi2 : entity work.handshake_addi_0(arch)
    port map(
      lhs => extsi8_outs,
      lhs_valid => extsi8_outs_valid,
      lhs_ready => extsi8_outs_ready,
      rhs => extsi16_outs,
      rhs_valid => extsi16_outs_valid,
      rhs_ready => extsi16_outs_ready,
      clk => clk,
      rst => rst,
      result => addi2_result,
      result_valid => addi2_result_valid,
      result_ready => addi2_result_ready
    );

  fork11 : entity work.handshake_fork_6(arch)
    port map(
      ins => addi2_result,
      ins_valid => addi2_result_valid,
      ins_ready => addi2_result_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork11_outs_0,
      outs(1) => fork11_outs_1,
      outs_valid(0) => fork11_outs_0_valid,
      outs_valid(1) => fork11_outs_1_valid,
      outs_ready(0) => fork11_outs_0_ready,
      outs_ready(1) => fork11_outs_1_ready
    );

  buffer191 : entity work.handshake_buffer_7(arch)
    port map(
      ins => fork11_outs_1,
      ins_valid => fork11_outs_1_valid,
      ins_ready => fork11_outs_1_ready,
      clk => clk,
      rst => rst,
      outs => buffer191_outs,
      outs_valid => buffer191_outs_valid,
      outs_ready => buffer191_outs_ready
    );

  buffer192 : entity work.handshake_buffer_7(arch)
    port map(
      ins => buffer191_outs,
      ins_valid => buffer191_outs_valid,
      ins_ready => buffer191_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer192_outs,
      outs_valid => buffer192_outs_valid,
      outs_ready => buffer192_outs_ready
    );

  buffer193 : entity work.handshake_buffer_7(arch)
    port map(
      ins => buffer192_outs,
      ins_valid => buffer192_outs_valid,
      ins_ready => buffer192_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer193_outs,
      outs_valid => buffer193_outs_valid,
      outs_ready => buffer193_outs_ready
    );

  buffer194 : entity work.handshake_buffer_7(arch)
    port map(
      ins => buffer193_outs,
      ins_valid => buffer193_outs_valid,
      ins_ready => buffer193_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer194_outs,
      outs_valid => buffer194_outs_valid,
      outs_ready => buffer194_outs_ready
    );

  buffer195 : entity work.handshake_buffer_7(arch)
    port map(
      ins => buffer194_outs,
      ins_valid => buffer194_outs_valid,
      ins_ready => buffer194_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer195_outs,
      outs_valid => buffer195_outs_valid,
      outs_ready => buffer195_outs_ready
    );

  trunci2 : entity work.handshake_trunci_1(arch)
    port map(
      ins => buffer195_outs,
      ins_valid => buffer195_outs_valid,
      ins_ready => buffer195_outs_ready,
      clk => clk,
      rst => rst,
      outs => trunci2_outs,
      outs_valid => trunci2_outs_valid,
      outs_ready => trunci2_outs_ready
    );

  buffer186 : entity work.handshake_buffer_7(arch)
    port map(
      ins => fork11_outs_0,
      ins_valid => fork11_outs_0_valid,
      ins_ready => fork11_outs_0_ready,
      clk => clk,
      rst => rst,
      outs => buffer186_outs,
      outs_valid => buffer186_outs_valid,
      outs_ready => buffer186_outs_ready
    );

  buffer187 : entity work.handshake_buffer_7(arch)
    port map(
      ins => buffer186_outs,
      ins_valid => buffer186_outs_valid,
      ins_ready => buffer186_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer187_outs,
      outs_valid => buffer187_outs_valid,
      outs_ready => buffer187_outs_ready
    );

  buffer188 : entity work.handshake_buffer_7(arch)
    port map(
      ins => buffer187_outs,
      ins_valid => buffer187_outs_valid,
      ins_ready => buffer187_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer188_outs,
      outs_valid => buffer188_outs_valid,
      outs_ready => buffer188_outs_ready
    );

  buffer189 : entity work.handshake_buffer_7(arch)
    port map(
      ins => buffer188_outs,
      ins_valid => buffer188_outs_valid,
      ins_ready => buffer188_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer189_outs,
      outs_valid => buffer189_outs_valid,
      outs_ready => buffer189_outs_ready
    );

  buffer190 : entity work.handshake_buffer_7(arch)
    port map(
      ins => buffer189_outs,
      ins_valid => buffer189_outs_valid,
      ins_ready => buffer189_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer190_outs,
      outs_valid => buffer190_outs_valid,
      outs_ready => buffer190_outs_ready
    );

  cmpi1 : entity work.handshake_cmpi_0(arch)
    port map(
      lhs => buffer190_outs,
      lhs_valid => buffer190_outs_valid,
      lhs_ready => buffer190_outs_ready,
      rhs => extsi15_outs,
      rhs_valid => extsi15_outs_valid,
      rhs_ready => extsi15_outs_ready,
      clk => clk,
      rst => rst,
      result => cmpi1_result,
      result_valid => cmpi1_result_valid,
      result_ready => cmpi1_result_ready
    );

  fork12 : entity work.handshake_fork_8(arch)
    port map(
      ins => cmpi1_result,
      ins_valid => cmpi1_result_valid,
      ins_ready => cmpi1_result_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork12_outs_0,
      outs(1) => fork12_outs_1,
      outs(2) => fork12_outs_2,
      outs(3) => fork12_outs_3,
      outs_valid(0) => fork12_outs_0_valid,
      outs_valid(1) => fork12_outs_1_valid,
      outs_valid(2) => fork12_outs_2_valid,
      outs_valid(3) => fork12_outs_3_valid,
      outs_ready(0) => fork12_outs_0_ready,
      outs_ready(1) => fork12_outs_1_ready,
      outs_ready(2) => fork12_outs_2_ready,
      outs_ready(3) => fork12_outs_3_ready
    );

  buffer0 : entity work.handshake_buffer_0(arch)
    port map(
      ins_valid => fork0_outs_0_valid,
      ins_ready => fork0_outs_0_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer0_outs_valid,
      outs_ready => buffer0_outs_ready
    );

  buffer1 : entity work.handshake_buffer_0(arch)
    port map(
      ins_valid => buffer0_outs_valid,
      ins_ready => buffer0_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer1_outs_valid,
      outs_ready => buffer1_outs_ready
    );

  buffer2 : entity work.handshake_buffer_0(arch)
    port map(
      ins_valid => buffer1_outs_valid,
      ins_ready => buffer1_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer2_outs_valid,
      outs_ready => buffer2_outs_ready
    );

  buffer3 : entity work.handshake_buffer_0(arch)
    port map(
      ins_valid => buffer2_outs_valid,
      ins_ready => buffer2_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer3_outs_valid,
      outs_ready => buffer3_outs_ready
    );

  buffer4 : entity work.handshake_buffer_0(arch)
    port map(
      ins_valid => buffer3_outs_valid,
      ins_ready => buffer3_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer4_outs_valid,
      outs_ready => buffer4_outs_ready
    );

end architecture;
