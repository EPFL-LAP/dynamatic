module xls_addf32(
  input wire clk,
  input wire rst,
  input wire [31:0] rhs,
  input wire rhs_valid,
  input wire [31:0] lhs,
  input wire lhs_valid,
  input wire result_ready,
  output wire [31:0] result,
  output wire result_valid,
  output wire rhs_ready,
  output wire lhs_ready
);
  function automatic [3:0] priority_sel_4b_2way (input reg [1:0] sel, input reg [3:0] case0, input reg [3:0] case1, input reg [3:0] default_value);
    begin
      casez (sel)
        2'b?1: begin
          priority_sel_4b_2way = case0;
        end
        2'b10: begin
          priority_sel_4b_2way = case1;
        end
        2'b00: begin
          priority_sel_4b_2way = default_value;
        end
        default: begin
          // Propagate X
          priority_sel_4b_2way = 4'dx;
        end
      endcase
    end
  endfunction
  function automatic [1:0] priority_sel_2b_2way (input reg [1:0] sel, input reg [1:0] case0, input reg [1:0] case1, input reg [1:0] default_value);
    begin
      casez (sel)
        2'b?1: begin
          priority_sel_2b_2way = case0;
        end
        2'b10: begin
          priority_sel_2b_2way = case1;
        end
        2'b00: begin
          priority_sel_2b_2way = default_value;
        end
        default: begin
          // Propagate X
          priority_sel_2b_2way = 2'dx;
        end
      endcase
    end
  endfunction
  function automatic priority_sel_1b_4way (input reg [3:0] sel, input reg case0, input reg case1, input reg case2, input reg case3, input reg default_value);
    begin
      casez (sel)
        4'b???1: begin
          priority_sel_1b_4way = case0;
        end
        4'b??10: begin
          priority_sel_1b_4way = case1;
        end
        4'b?100: begin
          priority_sel_1b_4way = case2;
        end
        4'b1000: begin
          priority_sel_1b_4way = case3;
        end
        4'b0000: begin
          priority_sel_1b_4way = default_value;
        end
        default: begin
          // Propagate X
          priority_sel_1b_4way = 1'dx;
        end
      endcase
    end
  endfunction
  function automatic priority_sel_1b_3way (input reg [2:0] sel, input reg case0, input reg case1, input reg case2, input reg default_value);
    begin
      casez (sel)
        3'b??1: begin
          priority_sel_1b_3way = case0;
        end
        3'b?10: begin
          priority_sel_1b_3way = case1;
        end
        3'b100: begin
          priority_sel_1b_3way = case2;
        end
        3'b000: begin
          priority_sel_1b_3way = default_value;
        end
        default: begin
          // Propagate X
          priority_sel_1b_3way = 1'dx;
        end
      endcase
    end
  endfunction
  function automatic [2:0] priority_sel_3b_2way (input reg [1:0] sel, input reg [2:0] case0, input reg [2:0] case1, input reg [2:0] default_value);
    begin
      casez (sel)
        2'b?1: begin
          priority_sel_3b_2way = case0;
        end
        2'b10: begin
          priority_sel_3b_2way = case1;
        end
        2'b00: begin
          priority_sel_3b_2way = default_value;
        end
        default: begin
          // Propagate X
          priority_sel_3b_2way = 3'dx;
        end
      endcase
    end
  endfunction
  function automatic [1:0] priority_sel_2b_4way (input reg [3:0] sel, input reg [1:0] case0, input reg [1:0] case1, input reg [1:0] case2, input reg [1:0] case3, input reg [1:0] default_value);
    begin
      casez (sel)
        4'b???1: begin
          priority_sel_2b_4way = case0;
        end
        4'b??10: begin
          priority_sel_2b_4way = case1;
        end
        4'b?100: begin
          priority_sel_2b_4way = case2;
        end
        4'b1000: begin
          priority_sel_2b_4way = case3;
        end
        4'b0000: begin
          priority_sel_2b_4way = default_value;
        end
        default: begin
          // Propagate X
          priority_sel_2b_4way = 2'dx;
        end
      endcase
    end
  endfunction
  function automatic priority_sel_1b_2way (input reg [1:0] sel, input reg case0, input reg case1, input reg default_value);
    begin
      casez (sel)
        2'b?1: begin
          priority_sel_1b_2way = case0;
        end
        2'b10: begin
          priority_sel_1b_2way = case1;
        end
        2'b00: begin
          priority_sel_1b_2way = default_value;
        end
        default: begin
          // Propagate X
          priority_sel_1b_2way = 1'dx;
        end
      endcase
    end
  endfunction
  wire [31:0] rhs_reg_init = {1'h0, 8'h00, 23'h00_0000};
  wire [31:0] lhs_reg_init = {1'h0, 8'h00, 23'h00_0000};
  wire [31:0] result_reg_init = {1'h0, 8'h00, 23'h00_0000};
  reg [7:0] p0_b_bexp__3;
  reg [7:0] p0_a_bexp__1;
  reg p0_bit_slice_20520;
  reg [22:0] p0_tuple_index_20521;
  reg [22:0] p0_tuple_index_20522;
  reg [7:0] p0_bit_slice_20523;
  reg p0_tuple_index_20524;
  reg p0_tuple_index_20525;
  reg [7:0] p1_a_bexp;
  reg p1_b_sign;
  reg p1_xor_20579;
  reg [24:0] p1_wide_x_squeezed;
  reg [24:0] p1_bit_slice_20581;
  reg [27:0] p1_shrl_20582;
  reg p1_sticky;
  reg p1_is_operand_inf;
  reg p1_and_20612;
  reg p1_is_result_nan;
  reg p1_not_20614;
  reg [7:0] p2_a_bexp;
  reg [27:0] p2_abs_fraction;
  reg p2_not_20660;
  reg p2_is_operand_inf;
  reg p2_is_result_nan;
  reg p2_result_sign;
  reg p2_not_20614;
  reg [7:0] p3_a_bexp;
  reg [27:0] p3_abs_fraction;
  reg p3_carry_bit;
  reg p3_and_20801;
  reg p3_and_20803;
  reg p3_nor_20809;
  reg p3_nor_20836;
  reg p3_and_20837;
  reg [2:0] p3_priority_sel_20838;
  reg [1:0] p3_priority_sel_20839;
  reg [2:0] p3_priority_sel_20840;
  reg p3_or_20841;
  reg p3_not_20660;
  reg p3_is_operand_inf;
  reg p3_is_result_nan;
  reg p3_result_sign__2;
  reg [7:0] p4_a_bexp;
  reg p4_and_20837;
  reg [3:0] p4_leading_zeroes__0_to_4;
  reg [2:0] p4_normal_chunk;
  reg [1:0] p4_half_way_chunk;
  reg [23:0] p4_bit_slice_20895;
  reg p4_not_20660;
  reg p4_is_operand_inf;
  reg p4_is_result_nan;
  reg p4_result_sign__2;
  reg p5_and_20837;
  reg [3:0] p5_leading_zeroes__0_to_4;
  reg [9:0] p5_concat_20935;
  reg p5_not_20660;
  reg p5_is_operand_inf;
  reg p5_is_result_nan;
  reg [22:0] p5_result_fraction;
  reg p5_result_sign__2;
  reg [8:0] p6_wide_exponent__2;
  reg p6_is_operand_inf;
  reg p6_is_result_nan;
  reg [22:0] p6_result_fraction;
  reg p6_result_sign__2;
  reg p7_is_result_nan;
  reg [22:0] p7_result_fraction__3;
  reg p7_result_sign__2;
  reg [7:0] p7_result_exponent__2;
  reg p0_valid;
  reg p1_valid;
  reg p2_valid;
  reg p3_valid;
  reg p4_valid;
  reg p5_valid;
  reg p6_valid;
  reg p7_valid;
  reg [31:0] rhs_reg;
  reg rhs_valid_reg;
  reg [31:0] lhs_reg;
  reg lhs_valid_reg;
  reg [31:0] result_reg;
  reg result_valid_reg;
  wire result_valid_inv;
  wire result_valid_load_en;
  wire result_load_en;
  wire p8_stage_done;
  wire p8_not_valid;
  wire p7_enable;
  wire p7_data_enable;
  wire p7_not_valid;
  wire p6_enable;
  wire p6_data_enable;
  wire p6_not_valid;
  wire p5_enable;
  wire p5_data_enable;
  wire p5_not_valid;
  wire p4_enable;
  wire p4_data_enable;
  wire p4_not_valid;
  wire p3_enable;
  wire p3_data_enable;
  wire p3_not_valid;
  wire [2:0] fraction_shift__3;
  wire p2_enable;
  wire [9:0] add_20962;
  wire [24:0] concat_20923;
  wire carry_bit;
  wire [24:0] addend_x__1_squeezed;
  wire [7:0] a_bexp;
  wire [7:0] incremented_sum__1;
  wire [7:0] MAX_EXPONENT;
  wire [22:0] a_fraction;
  wire [7:0] b_bexp;
  wire [7:0] MAX_EXPONENT__1;
  wire [22:0] b_fraction;
  wire p2_data_enable;
  wire p2_not_valid;
  wire [9:0] wide_exponent;
  wire do_round_up;
  wire [24:0] add_20926;
  wire [3:0] leading_zeroes__0_to_4;
  wire nor_20708;
  wire nor_20709;
  wire nor_20711;
  wire nor_20712;
  wire nor_20717;
  wire nor_20718;
  wire nor_20723;
  wire nor_20726;
  wire nor_20727;
  wire nor_20728;
  wire nor_20734;
  wire [7:0] a_bexpbs_difference__1;
  wire eq_20592;
  wire eq_20593;
  wire eq_20594;
  wire eq_20595;
  wire p1_enable;
  wire and_reduce_20989;
  wire [9:0] wide_exponent__1;
  wire [24:0] rounded_fraction_squeezed_portion_3_width_25;
  wire [4:0] leading_zeroes;
  wire nor_20735;
  wire and_20736;
  wire and_20738;
  wire nor_20743;
  wire and_20744;
  wire nor_20747;
  wire and_20751;
  wire nor_20752;
  wire and_20756;
  wire nor_20758;
  wire [25:0] add_20644;
  wire [23:0] fraction_x;
  wire a_sign;
  wire b_sign;
  wire [7:0] b_bexp__3;
  wire p1_data_enable;
  wire p1_not_valid;
  wire rounding_carry;
  wire [2:0] fraction_shift__2;
  wire [2:0] fraction_shift__4;
  wire [28:0] cancel_fraction;
  wire and_20765;
  wire and_20783;
  wire [23:0] fraction_x__1;
  wire [2:0] addend_x__1_squeezed_const_lsb_bits__1;
  wire [23:0] fraction_y;
  wire [23:0] sign_ext_20564;
  wire [27:0] add_20583;
  wire [7:0] a_bexp__1;
  wire p0_enable;
  wire p0_all_active_inputs_valid;
  wire [27:0] rounded_fraction;
  wire [2:0] fraction_shift__1;
  wire [26:0] cancel_fraction__1;
  wire [26:0] carry_fraction__1;
  wire and_20801;
  wire and_20803;
  wire nor_20809;
  wire and_20810;
  wire [1:0] priority_sel_20817;
  wire [27:0] concat_20649;
  wire fraction_is_zero;
  wire [27:0] wide_x;
  wire [23:0] fraction_y__1;
  wire [2:0] addend_x__1_squeezed_const_lsb_bits;
  wire has_pos_inf;
  wire has_neg_inf;
  wire p0_data_enable;
  wire rhs_valid_inv;
  wire lhs_valid_inv;
  wire [22:0] FRACTION_HIGH_BIT;
  wire [7:0] MAX_EXPONENT__2;
  wire [8:0] add_20934;
  wire [27:0] shrl_20940;
  wire [26:0] shifted_fraction;
  wire result_sign__1;
  wire [27:0] neg_20575;
  wire [27:0] wide_y;
  wire [8:0] sum__1;
  wire rhs_valid_load_en;
  wire lhs_valid_load_en;
  wire [22:0] result_fraction__4;
  wire [22:0] result_fraction__3;
  wire [7:0] result_exponent__2;
  wire [8:0] wide_exponent__2;
  wire [9:0] concat_20935;
  wire [22:0] result_fraction;
  wire [2:0] normal_chunk;
  wire [1:0] half_way_chunk;
  wire [23:0] bit_slice_20895;
  wire nor_20836;
  wire and_20837;
  wire [2:0] priority_sel_20838;
  wire [1:0] priority_sel_20839;
  wire [2:0] priority_sel_20840;
  wire or_20841;
  wire result_sign__2;
  wire [27:0] abs_fraction;
  wire not_20660;
  wire result_sign;
  wire xor_20579;
  wire [24:0] wide_x_squeezed;
  wire [24:0] bit_slice_20581;
  wire [27:0] shrl_20582;
  wire sticky;
  wire is_operand_inf;
  wire and_20612;
  wire is_result_nan;
  wire not_20614;
  wire bit_slice_20520;
  wire [22:0] tuple_index_20521;
  wire [22:0] tuple_index_20522;
  wire [7:0] bit_slice_20523;
  wire tuple_index_20524;
  wire tuple_index_20525;
  wire rhs_load_en;
  wire lhs_load_en;
  wire [31:0] sum;
  assign result_valid_inv = ~result_valid_reg;
  assign result_valid_load_en = result_ready | result_valid_inv;
  assign result_load_en = p7_valid & result_valid_load_en;
  assign p8_stage_done = p7_valid & result_load_en;
  assign p8_not_valid = ~p7_valid;
  assign p7_enable = p8_stage_done | p8_not_valid;
  assign p7_data_enable = p7_enable & p6_valid;
  assign p7_not_valid = ~p6_valid;
  assign p6_enable = p7_data_enable | p7_not_valid;
  assign p6_data_enable = p6_enable & p5_valid;
  assign p6_not_valid = ~p5_valid;
  assign p5_enable = p6_data_enable | p6_not_valid;
  assign p5_data_enable = p5_enable & p4_valid;
  assign p5_not_valid = ~p4_valid;
  assign p4_enable = p5_data_enable | p5_not_valid;
  assign p4_data_enable = p4_enable & p3_valid;
  assign p4_not_valid = ~p3_valid;
  assign p3_enable = p4_data_enable | p4_not_valid;
  assign p3_data_enable = p3_enable & p2_valid;
  assign p3_not_valid = ~p2_valid;
  assign fraction_shift__3 = 3'h4;
  assign p2_enable = p3_data_enable | p3_not_valid;
  assign add_20962 = p5_concat_20935 + 10'h001;
  assign concat_20923 = {1'h0, p4_bit_slice_20895};
  assign carry_bit = p2_abs_fraction[27];
  assign addend_x__1_squeezed = p1_xor_20579 ? p1_bit_slice_20581 : p1_wide_x_squeezed;
  assign a_bexp = p0_bit_slice_20520 ? p0_a_bexp__1 : p0_b_bexp__3;
  assign incremented_sum__1 = p0_bit_slice_20523 + 8'h01;
  assign MAX_EXPONENT = 8'hff;
  assign a_fraction = p0_bit_slice_20520 ? p0_tuple_index_20522 : p0_tuple_index_20521;
  assign b_bexp = p0_bit_slice_20520 ? p0_b_bexp__3 : p0_a_bexp__1;
  assign MAX_EXPONENT__1 = 8'hff;
  assign b_fraction = p0_bit_slice_20520 ? p0_tuple_index_20521 : p0_tuple_index_20522;
  assign p2_data_enable = p2_enable & p1_valid;
  assign p2_not_valid = ~p1_valid;
  assign wide_exponent = add_20962 - {5'h00, p5_and_20837, p5_leading_zeroes__0_to_4};
  assign do_round_up = p4_normal_chunk > fraction_shift__3 | p4_half_way_chunk == 2'h3;
  assign add_20926 = concat_20923 + 25'h000_0001;
  assign leading_zeroes__0_to_4 = priority_sel_4b_2way({p3_nor_20836, p3_and_20837}, {p3_and_20803, p3_priority_sel_20838}, {1'h1, p3_nor_20809, p3_priority_sel_20839}, {p3_and_20801, p3_priority_sel_20840});
  assign nor_20708 = ~(p2_abs_fraction[11] | p2_abs_fraction[10]);
  assign nor_20709 = ~(p2_abs_fraction[9] | p2_abs_fraction[8]);
  assign nor_20711 = ~(p2_abs_fraction[1] | p2_abs_fraction[0]);
  assign nor_20712 = ~(p2_abs_fraction[3] | p2_abs_fraction[2]);
  assign nor_20717 = ~(p2_abs_fraction[5] | p2_abs_fraction[4]);
  assign nor_20718 = ~(p2_abs_fraction[7] | p2_abs_fraction[6]);
  assign nor_20723 = ~(p2_abs_fraction[17] | p2_abs_fraction[16]);
  assign nor_20726 = ~(p2_abs_fraction[13] | p2_abs_fraction[12]);
  assign nor_20727 = ~(carry_bit | p2_abs_fraction[26]);
  assign nor_20728 = ~(p2_abs_fraction[25] | p2_abs_fraction[24]);
  assign nor_20734 = ~(p2_abs_fraction[21] | p2_abs_fraction[20]);
  assign a_bexpbs_difference__1 = p0_bit_slice_20520 ? incremented_sum__1 : ~p0_bit_slice_20523;
  assign eq_20592 = a_bexp == MAX_EXPONENT;
  assign eq_20593 = a_fraction == 23'h00_0000;
  assign eq_20594 = b_bexp == MAX_EXPONENT__1;
  assign eq_20595 = b_fraction == 23'h00_0000;
  assign p1_enable = p2_data_enable | p2_not_valid;
  assign and_reduce_20989 = &p6_wide_exponent__2[7:0];
  assign wide_exponent__1 = wide_exponent & {10{p5_not_20660}};
  assign rounded_fraction_squeezed_portion_3_width_25 = do_round_up ? add_20926 : concat_20923;
  assign leading_zeroes = {p3_and_20837, leading_zeroes__0_to_4};
  assign nor_20735 = ~(p2_abs_fraction[23] | p2_abs_fraction[22]);
  assign and_20736 = nor_20708 & nor_20709;
  assign and_20738 = nor_20712 & nor_20711;
  assign nor_20743 = ~(p2_abs_fraction[7] | p2_abs_fraction[6] | nor_20717);
  assign and_20744 = nor_20718 & nor_20717;
  assign nor_20747 = ~(p2_abs_fraction[11] | ~p2_abs_fraction[10]);
  assign and_20751 = ~(p2_abs_fraction[19] | p2_abs_fraction[18]) & nor_20723;
  assign nor_20752 = ~(p2_abs_fraction[15] | p2_abs_fraction[14]);
  assign and_20756 = nor_20727 & nor_20728;
  assign nor_20758 = ~(carry_bit | ~p2_abs_fraction[26]);
  assign add_20644 = {{1{addend_x__1_squeezed[24]}}, addend_x__1_squeezed} + {1'h0, p1_shrl_20582[27:3]};
  assign fraction_x = {1'h1, a_fraction};
  assign a_sign = p0_bit_slice_20520 ? p0_tuple_index_20525 : p0_tuple_index_20524;
  assign b_sign = p0_bit_slice_20520 ? p0_tuple_index_20524 : p0_tuple_index_20525;
  assign b_bexp__3 = rhs_reg[30:23];
  assign p1_data_enable = p1_enable & p0_valid;
  assign p1_not_valid = ~p0_valid;
  assign rounding_carry = rounded_fraction_squeezed_portion_3_width_25[24];
  assign fraction_shift__2 = 3'h3;
  assign fraction_shift__4 = 3'h4;
  assign cancel_fraction = leading_zeroes >= 5'h1d ? 29'h0000_0000 : {1'h0, p3_abs_fraction} << leading_zeroes;
  assign and_20765 = nor_20735 & nor_20734;
  assign and_20783 = nor_20752 & nor_20726;
  assign fraction_x__1 = fraction_x & {24{a_bexp != 8'h00}};
  assign addend_x__1_squeezed_const_lsb_bits__1 = 3'h0;
  assign fraction_y = {1'h1, b_fraction};
  assign sign_ext_20564 = {24{b_bexp != 8'h00}};
  assign add_20583 = (a_bexpbs_difference__1 >= 8'h1c ? 28'h000_0000 : 28'h000_0001 << a_bexpbs_difference__1) + 28'hfff_ffff;
  assign a_bexp__1 = lhs_reg[30:23];
  assign p0_enable = p1_data_enable | p1_not_valid;
  assign p0_all_active_inputs_valid = rhs_valid_reg & lhs_valid_reg;
  assign rounded_fraction = {rounded_fraction_squeezed_portion_3_width_25, p4_normal_chunk};
  assign fraction_shift__1 = rounding_carry ? fraction_shift__4 : fraction_shift__2;
  assign cancel_fraction__1 = cancel_fraction[27:1];
  assign carry_fraction__1 = {p3_abs_fraction[27:2], p3_or_20841};
  assign and_20801 = and_20756 & and_20765;
  assign and_20803 = and_20736 & and_20744;
  assign nor_20809 = ~(~and_20751 | and_20783);
  assign and_20810 = and_20751 & and_20783;
  assign priority_sel_20817 = priority_sel_2b_2way({~(carry_bit | p2_abs_fraction[26] | nor_20728), and_20756}, {nor_20758, 1'h0}, {1'h1, ~(p2_abs_fraction[25] | ~p2_abs_fraction[24])}, {nor_20727, nor_20758});
  assign concat_20649 = {add_20644[24:0], p1_shrl_20582[2:1], p1_shrl_20582[0] | p1_sticky};
  assign fraction_is_zero = add_20644 == 26'h000_0000 & ~(p1_shrl_20582[1] | p1_shrl_20582[2]) & ~(p1_shrl_20582[0] | p1_sticky);
  assign wide_x = {1'h0, fraction_x__1, addend_x__1_squeezed_const_lsb_bits__1};
  assign fraction_y__1 = fraction_y & sign_ext_20564;
  assign addend_x__1_squeezed_const_lsb_bits = 3'h0;
  assign has_pos_inf = ~(~eq_20592 | ~eq_20593 | a_sign) | ~(~eq_20594 | ~eq_20595 | b_sign);
  assign has_neg_inf = eq_20592 & eq_20593 & a_sign | eq_20594 & eq_20595 & b_sign;
  assign p0_data_enable = p0_enable & p0_all_active_inputs_valid;
  assign rhs_valid_inv = ~rhs_valid_reg;
  assign lhs_valid_inv = ~lhs_valid_reg;
  assign FRACTION_HIGH_BIT = 23'h40_0000;
  assign MAX_EXPONENT__2 = 8'hff;
  assign add_20934 = {1'h0, p4_a_bexp} + {8'h00, rounding_carry};
  assign shrl_20940 = rounded_fraction >> fraction_shift__1;
  assign shifted_fraction = p3_carry_bit ? carry_fraction__1 : cancel_fraction__1;
  assign result_sign__1 = p2_is_operand_inf ? p2_not_20614 : p2_result_sign;
  assign neg_20575 = -wide_x;
  assign wide_y = {1'h0, fraction_y__1, addend_x__1_squeezed_const_lsb_bits};
  assign sum__1 = {1'h0, a_bexp__1} + {1'h0, ~b_bexp__3};
  assign rhs_valid_load_en = p0_data_enable | rhs_valid_inv;
  assign lhs_valid_load_en = p0_data_enable | lhs_valid_inv;
  assign result_fraction__4 = p7_is_result_nan ? FRACTION_HIGH_BIT : p7_result_fraction__3;
  assign result_fraction__3 = p6_result_fraction & {23{~(p6_is_operand_inf | p6_wide_exponent__2[8] | and_reduce_20989 | ~((|p6_wide_exponent__2[8:1]) | p6_wide_exponent__2[0]))}};
  assign result_exponent__2 = p6_is_result_nan | p6_is_operand_inf | p6_wide_exponent__2[8] | and_reduce_20989 ? MAX_EXPONENT__2 : p6_wide_exponent__2[7:0];
  assign wide_exponent__2 = wide_exponent__1[8:0] & {9{~wide_exponent__1[9]}};
  assign concat_20935 = {1'h0, add_20934};
  assign result_fraction = shrl_20940[22:0];
  assign normal_chunk = shifted_fraction[2:0];
  assign half_way_chunk = shifted_fraction[3:2];
  assign bit_slice_20895 = shifted_fraction[26:3];
  assign nor_20836 = ~(~and_20801 | and_20810);
  assign and_20837 = and_20801 & and_20810;
  assign priority_sel_20838 = priority_sel_3b_2way({~(~and_20736 | and_20744), and_20803}, {and_20738, priority_sel_2b_2way({~(p2_abs_fraction[3] | p2_abs_fraction[2] | nor_20711), and_20738}, 2'h0, {1'h1, ~(p2_abs_fraction[1] | ~p2_abs_fraction[0])}, {nor_20712, ~(p2_abs_fraction[3] | ~p2_abs_fraction[2])})}, {1'h1, nor_20743, priority_sel_1b_4way({~(p2_abs_fraction[7] | ~p2_abs_fraction[6]), nor_20718, nor_20743, and_20744}, 1'h0, ~(p2_abs_fraction[5] | ~p2_abs_fraction[4]), 1'h0, 1'h1, 1'h0)}, {and_20736, priority_sel_2b_2way({~(p2_abs_fraction[11] | p2_abs_fraction[10] | nor_20709), and_20736}, {nor_20747, 1'h0}, {1'h1, ~(p2_abs_fraction[9] | ~p2_abs_fraction[8])}, {nor_20708, nor_20747})});
  assign priority_sel_20839 = priority_sel_2b_4way({~(p2_abs_fraction[19] | p2_abs_fraction[18] | nor_20723), and_20751, nor_20809, and_20810}, 2'h0, {nor_20752, priority_sel_1b_3way({~(p2_abs_fraction[15] | ~p2_abs_fraction[14]), nor_20752, ~(p2_abs_fraction[15] | p2_abs_fraction[14] | nor_20726)}, ~(p2_abs_fraction[13] | ~p2_abs_fraction[12]), 1'h0, 1'h1, 1'h0)}, 2'h0, {1'h1, ~(p2_abs_fraction[17] | ~p2_abs_fraction[16])}, {1'h0, ~(p2_abs_fraction[19] | ~p2_abs_fraction[18])});
  assign priority_sel_20840 = priority_sel_3b_2way({~(~and_20756 | and_20765), and_20801}, {priority_sel_20817, 1'h0}, {1'h1, nor_20735, priority_sel_1b_3way({~(p2_abs_fraction[23] | ~p2_abs_fraction[22]), nor_20735, ~(p2_abs_fraction[23] | p2_abs_fraction[22] | nor_20734)}, ~(p2_abs_fraction[21] | ~p2_abs_fraction[20]), 1'h0, 1'h1, 1'h0)}, {and_20756, priority_sel_20817});
  assign or_20841 = p2_abs_fraction[1] | p2_abs_fraction[0];
  assign result_sign__2 = ~p2_is_result_nan & result_sign__1;
  assign abs_fraction = add_20644[25] ? -concat_20649 : concat_20649;
  assign not_20660 = ~fraction_is_zero;
  assign result_sign = priority_sel_1b_2way({add_20644[25], fraction_is_zero}, p1_and_20612, ~p1_b_sign, p1_b_sign);
  assign xor_20579 = a_sign ^ b_sign;
  assign wide_x_squeezed = {1'h0, fraction_x__1};
  assign bit_slice_20581 = neg_20575[27:3];
  assign shrl_20582 = a_bexpbs_difference__1 >= 8'h1c ? 28'h000_0000 : wide_y >> a_bexpbs_difference__1;
  assign sticky = (fraction_y & sign_ext_20564 & add_20583[26:3]) != 24'h00_0000;
  assign is_operand_inf = eq_20592 & eq_20593 | eq_20594 & eq_20595;
  assign and_20612 = a_sign & b_sign;
  assign is_result_nan = ~(~eq_20592 | eq_20593) | ~(~eq_20594 | eq_20595) | has_pos_inf & has_neg_inf;
  assign not_20614 = ~has_pos_inf;
  assign bit_slice_20520 = sum__1[8];
  assign tuple_index_20521 = rhs_reg[22:0];
  assign tuple_index_20522 = lhs_reg[22:0];
  assign bit_slice_20523 = sum__1[7:0];
  assign tuple_index_20524 = rhs_reg[31:31];
  assign tuple_index_20525 = lhs_reg[31:31];
  assign rhs_load_en = rhs_valid & rhs_valid_load_en;
  assign lhs_load_en = lhs_valid & lhs_valid_load_en;
  assign sum = {p7_result_sign__2, p7_result_exponent__2, result_fraction__4};
  always @ (posedge clk) begin
    if (rst) begin
      p0_b_bexp__3 <= 8'h00;
      p0_a_bexp__1 <= 8'h00;
      p0_bit_slice_20520 <= 1'h0;
      p0_tuple_index_20521 <= 23'h00_0000;
      p0_tuple_index_20522 <= 23'h00_0000;
      p0_bit_slice_20523 <= 8'h00;
      p0_tuple_index_20524 <= 1'h0;
      p0_tuple_index_20525 <= 1'h0;
      p1_a_bexp <= 8'h00;
      p1_b_sign <= 1'h0;
      p1_xor_20579 <= 1'h0;
      p1_wide_x_squeezed <= 25'h000_0000;
      p1_bit_slice_20581 <= 25'h000_0000;
      p1_shrl_20582 <= 28'h000_0000;
      p1_sticky <= 1'h0;
      p1_is_operand_inf <= 1'h0;
      p1_and_20612 <= 1'h0;
      p1_is_result_nan <= 1'h0;
      p1_not_20614 <= 1'h0;
      p2_a_bexp <= 8'h00;
      p2_abs_fraction <= 28'h000_0000;
      p2_not_20660 <= 1'h0;
      p2_is_operand_inf <= 1'h0;
      p2_is_result_nan <= 1'h0;
      p2_result_sign <= 1'h0;
      p2_not_20614 <= 1'h0;
      p3_a_bexp <= 8'h00;
      p3_abs_fraction <= 28'h000_0000;
      p3_carry_bit <= 1'h0;
      p3_and_20801 <= 1'h0;
      p3_and_20803 <= 1'h0;
      p3_nor_20809 <= 1'h0;
      p3_nor_20836 <= 1'h0;
      p3_and_20837 <= 1'h0;
      p3_priority_sel_20838 <= 3'h0;
      p3_priority_sel_20839 <= 2'h0;
      p3_priority_sel_20840 <= 3'h0;
      p3_or_20841 <= 1'h0;
      p3_not_20660 <= 1'h0;
      p3_is_operand_inf <= 1'h0;
      p3_is_result_nan <= 1'h0;
      p3_result_sign__2 <= 1'h0;
      p4_a_bexp <= 8'h00;
      p4_and_20837 <= 1'h0;
      p4_leading_zeroes__0_to_4 <= 4'h0;
      p4_normal_chunk <= 3'h0;
      p4_half_way_chunk <= 2'h0;
      p4_bit_slice_20895 <= 24'h00_0000;
      p4_not_20660 <= 1'h0;
      p4_is_operand_inf <= 1'h0;
      p4_is_result_nan <= 1'h0;
      p4_result_sign__2 <= 1'h0;
      p5_and_20837 <= 1'h0;
      p5_leading_zeroes__0_to_4 <= 4'h0;
      p5_concat_20935 <= 10'h000;
      p5_not_20660 <= 1'h0;
      p5_is_operand_inf <= 1'h0;
      p5_is_result_nan <= 1'h0;
      p5_result_fraction <= 23'h00_0000;
      p5_result_sign__2 <= 1'h0;
      p6_wide_exponent__2 <= 9'h000;
      p6_is_operand_inf <= 1'h0;
      p6_is_result_nan <= 1'h0;
      p6_result_fraction <= 23'h00_0000;
      p6_result_sign__2 <= 1'h0;
      p7_is_result_nan <= 1'h0;
      p7_result_fraction__3 <= 23'h00_0000;
      p7_result_sign__2 <= 1'h0;
      p7_result_exponent__2 <= 8'h00;
      p0_valid <= 1'h0;
      p1_valid <= 1'h0;
      p2_valid <= 1'h0;
      p3_valid <= 1'h0;
      p4_valid <= 1'h0;
      p5_valid <= 1'h0;
      p6_valid <= 1'h0;
      p7_valid <= 1'h0;
      rhs_reg <= rhs_reg_init;
      rhs_valid_reg <= 1'h0;
      lhs_reg <= lhs_reg_init;
      lhs_valid_reg <= 1'h0;
      result_reg <= result_reg_init;
      result_valid_reg <= 1'h0;
    end else begin
      p0_b_bexp__3 <= p0_data_enable ? b_bexp__3 : p0_b_bexp__3;
      p0_a_bexp__1 <= p0_data_enable ? a_bexp__1 : p0_a_bexp__1;
      p0_bit_slice_20520 <= p0_data_enable ? bit_slice_20520 : p0_bit_slice_20520;
      p0_tuple_index_20521 <= p0_data_enable ? tuple_index_20521 : p0_tuple_index_20521;
      p0_tuple_index_20522 <= p0_data_enable ? tuple_index_20522 : p0_tuple_index_20522;
      p0_bit_slice_20523 <= p0_data_enable ? bit_slice_20523 : p0_bit_slice_20523;
      p0_tuple_index_20524 <= p0_data_enable ? tuple_index_20524 : p0_tuple_index_20524;
      p0_tuple_index_20525 <= p0_data_enable ? tuple_index_20525 : p0_tuple_index_20525;
      p1_a_bexp <= p1_data_enable ? a_bexp : p1_a_bexp;
      p1_b_sign <= p1_data_enable ? b_sign : p1_b_sign;
      p1_xor_20579 <= p1_data_enable ? xor_20579 : p1_xor_20579;
      p1_wide_x_squeezed <= p1_data_enable ? wide_x_squeezed : p1_wide_x_squeezed;
      p1_bit_slice_20581 <= p1_data_enable ? bit_slice_20581 : p1_bit_slice_20581;
      p1_shrl_20582 <= p1_data_enable ? shrl_20582 : p1_shrl_20582;
      p1_sticky <= p1_data_enable ? sticky : p1_sticky;
      p1_is_operand_inf <= p1_data_enable ? is_operand_inf : p1_is_operand_inf;
      p1_and_20612 <= p1_data_enable ? and_20612 : p1_and_20612;
      p1_is_result_nan <= p1_data_enable ? is_result_nan : p1_is_result_nan;
      p1_not_20614 <= p1_data_enable ? not_20614 : p1_not_20614;
      p2_a_bexp <= p2_data_enable ? p1_a_bexp : p2_a_bexp;
      p2_abs_fraction <= p2_data_enable ? abs_fraction : p2_abs_fraction;
      p2_not_20660 <= p2_data_enable ? not_20660 : p2_not_20660;
      p2_is_operand_inf <= p2_data_enable ? p1_is_operand_inf : p2_is_operand_inf;
      p2_is_result_nan <= p2_data_enable ? p1_is_result_nan : p2_is_result_nan;
      p2_result_sign <= p2_data_enable ? result_sign : p2_result_sign;
      p2_not_20614 <= p2_data_enable ? p1_not_20614 : p2_not_20614;
      p3_a_bexp <= p3_data_enable ? p2_a_bexp : p3_a_bexp;
      p3_abs_fraction <= p3_data_enable ? p2_abs_fraction : p3_abs_fraction;
      p3_carry_bit <= p3_data_enable ? carry_bit : p3_carry_bit;
      p3_and_20801 <= p3_data_enable ? and_20801 : p3_and_20801;
      p3_and_20803 <= p3_data_enable ? and_20803 : p3_and_20803;
      p3_nor_20809 <= p3_data_enable ? nor_20809 : p3_nor_20809;
      p3_nor_20836 <= p3_data_enable ? nor_20836 : p3_nor_20836;
      p3_and_20837 <= p3_data_enable ? and_20837 : p3_and_20837;
      p3_priority_sel_20838 <= p3_data_enable ? priority_sel_20838 : p3_priority_sel_20838;
      p3_priority_sel_20839 <= p3_data_enable ? priority_sel_20839 : p3_priority_sel_20839;
      p3_priority_sel_20840 <= p3_data_enable ? priority_sel_20840 : p3_priority_sel_20840;
      p3_or_20841 <= p3_data_enable ? or_20841 : p3_or_20841;
      p3_not_20660 <= p3_data_enable ? p2_not_20660 : p3_not_20660;
      p3_is_operand_inf <= p3_data_enable ? p2_is_operand_inf : p3_is_operand_inf;
      p3_is_result_nan <= p3_data_enable ? p2_is_result_nan : p3_is_result_nan;
      p3_result_sign__2 <= p3_data_enable ? result_sign__2 : p3_result_sign__2;
      p4_a_bexp <= p4_data_enable ? p3_a_bexp : p4_a_bexp;
      p4_and_20837 <= p4_data_enable ? p3_and_20837 : p4_and_20837;
      p4_leading_zeroes__0_to_4 <= p4_data_enable ? leading_zeroes__0_to_4 : p4_leading_zeroes__0_to_4;
      p4_normal_chunk <= p4_data_enable ? normal_chunk : p4_normal_chunk;
      p4_half_way_chunk <= p4_data_enable ? half_way_chunk : p4_half_way_chunk;
      p4_bit_slice_20895 <= p4_data_enable ? bit_slice_20895 : p4_bit_slice_20895;
      p4_not_20660 <= p4_data_enable ? p3_not_20660 : p4_not_20660;
      p4_is_operand_inf <= p4_data_enable ? p3_is_operand_inf : p4_is_operand_inf;
      p4_is_result_nan <= p4_data_enable ? p3_is_result_nan : p4_is_result_nan;
      p4_result_sign__2 <= p4_data_enable ? p3_result_sign__2 : p4_result_sign__2;
      p5_and_20837 <= p5_data_enable ? p4_and_20837 : p5_and_20837;
      p5_leading_zeroes__0_to_4 <= p5_data_enable ? p4_leading_zeroes__0_to_4 : p5_leading_zeroes__0_to_4;
      p5_concat_20935 <= p5_data_enable ? concat_20935 : p5_concat_20935;
      p5_not_20660 <= p5_data_enable ? p4_not_20660 : p5_not_20660;
      p5_is_operand_inf <= p5_data_enable ? p4_is_operand_inf : p5_is_operand_inf;
      p5_is_result_nan <= p5_data_enable ? p4_is_result_nan : p5_is_result_nan;
      p5_result_fraction <= p5_data_enable ? result_fraction : p5_result_fraction;
      p5_result_sign__2 <= p5_data_enable ? p4_result_sign__2 : p5_result_sign__2;
      p6_wide_exponent__2 <= p6_data_enable ? wide_exponent__2 : p6_wide_exponent__2;
      p6_is_operand_inf <= p6_data_enable ? p5_is_operand_inf : p6_is_operand_inf;
      p6_is_result_nan <= p6_data_enable ? p5_is_result_nan : p6_is_result_nan;
      p6_result_fraction <= p6_data_enable ? p5_result_fraction : p6_result_fraction;
      p6_result_sign__2 <= p6_data_enable ? p5_result_sign__2 : p6_result_sign__2;
      p7_is_result_nan <= p7_data_enable ? p6_is_result_nan : p7_is_result_nan;
      p7_result_fraction__3 <= p7_data_enable ? result_fraction__3 : p7_result_fraction__3;
      p7_result_sign__2 <= p7_data_enable ? p6_result_sign__2 : p7_result_sign__2;
      p7_result_exponent__2 <= p7_data_enable ? result_exponent__2 : p7_result_exponent__2;
      p0_valid <= p0_enable ? p0_all_active_inputs_valid : p0_valid;
      p1_valid <= p1_enable ? p0_valid : p1_valid;
      p2_valid <= p2_enable ? p1_valid : p2_valid;
      p3_valid <= p3_enable ? p2_valid : p3_valid;
      p4_valid <= p4_enable ? p3_valid : p4_valid;
      p5_valid <= p5_enable ? p4_valid : p5_valid;
      p6_valid <= p6_enable ? p5_valid : p6_valid;
      p7_valid <= p7_enable ? p6_valid : p7_valid;
      rhs_reg <= rhs_load_en ? rhs : rhs_reg;
      rhs_valid_reg <= rhs_valid_load_en ? rhs_valid : rhs_valid_reg;
      lhs_reg <= lhs_load_en ? lhs : lhs_reg;
      lhs_valid_reg <= lhs_valid_load_en ? lhs_valid : lhs_valid_reg;
      result_reg <= result_load_en ? sum : result_reg;
      result_valid_reg <= result_valid_load_en ? p7_valid : result_valid_reg;
    end
  end
  assign result = result_reg;
  assign result_valid = result_valid_reg;
  assign rhs_ready = rhs_load_en;
  assign lhs_ready = lhs_load_en;
endmodule
module xls_cmpf32_OEQ(
  input wire clk,
  input wire rst,
  input wire [31:0] lhs,
  input wire lhs_valid,
  input wire [31:0] rhs,
  input wire rhs_valid,
  input wire result_ready,
  output wire result,
  output wire result_valid,
  output wire lhs_ready,
  output wire rhs_ready
);
  wire [31:0] lhs_reg_init = {1'h0, 8'h00, 23'h00_0000};
  wire [31:0] rhs_reg_init = {1'h0, 8'h00, 23'h00_0000};
  reg [31:0] lhs_reg;
  reg lhs_valid_reg;
  reg [31:0] rhs_reg;
  reg rhs_valid_reg;
  reg result_reg;
  reg result_valid_reg;
  wire result_valid_inv;
  wire p0_all_active_inputs_valid;
  wire result_valid_load_en;
  wire [7:0] a_bexp__4;
  wire [22:0] a_fraction__1;
  wire [7:0] b_bexp__1;
  wire [22:0] b_fraction__1;
  wire a_sign__1;
  wire b_sign;
  wire result_load_en;
  wire p0_stage_done;
  wire lhs_valid_inv;
  wire rhs_valid_inv;
  wire lhs_valid_load_en;
  wire rhs_valid_load_en;
  wire lhs_load_en;
  wire rhs_load_en;
  wire sum;
  assign result_valid_inv = ~result_valid_reg;
  assign p0_all_active_inputs_valid = lhs_valid_reg & rhs_valid_reg;
  assign result_valid_load_en = result_ready | result_valid_inv;
  assign a_bexp__4 = lhs_reg[30:23];
  assign a_fraction__1 = lhs_reg[22:0];
  assign b_bexp__1 = rhs_reg[30:23];
  assign b_fraction__1 = rhs_reg[22:0];
  assign a_sign__1 = lhs_reg[31:31];
  assign b_sign = rhs_reg[31:31];
  assign result_load_en = p0_all_active_inputs_valid & result_valid_load_en;
  assign p0_stage_done = p0_all_active_inputs_valid & result_load_en;
  assign lhs_valid_inv = ~lhs_valid_reg;
  assign rhs_valid_inv = ~rhs_valid_reg;
  assign lhs_valid_load_en = p0_stage_done | lhs_valid_inv;
  assign rhs_valid_load_en = p0_stage_done | rhs_valid_inv;
  assign lhs_load_en = lhs_valid & lhs_valid_load_en;
  assign rhs_load_en = rhs_valid & rhs_valid_load_en;
  assign sum = ~(a_bexp__4 == 8'hff & a_fraction__1 != 23'h00_0000 | b_bexp__1 == 8'hff & b_fraction__1 != 23'h00_0000) & (a_sign__1 == b_sign & a_bexp__4 == b_bexp__1 & a_fraction__1 == b_fraction__1 | a_bexp__4 == 8'h00 & b_bexp__1 == 8'h00);
  always @ (posedge clk) begin
    if (rst) begin
      lhs_reg <= lhs_reg_init;
      lhs_valid_reg <= 1'h0;
      rhs_reg <= rhs_reg_init;
      rhs_valid_reg <= 1'h0;
      result_reg <= 1'h0;
      result_valid_reg <= 1'h0;
    end else begin
      lhs_reg <= lhs_load_en ? lhs : lhs_reg;
      lhs_valid_reg <= lhs_valid_load_en ? lhs_valid : lhs_valid_reg;
      rhs_reg <= rhs_load_en ? rhs : rhs_reg;
      rhs_valid_reg <= rhs_valid_load_en ? rhs_valid : rhs_valid_reg;
      result_reg <= result_load_en ? sum : result_reg;
      result_valid_reg <= result_valid_load_en ? p0_all_active_inputs_valid : result_valid_reg;
    end
  end
  assign result = result_reg;
  assign result_valid = result_valid_reg;
  assign lhs_ready = lhs_load_en;
  assign rhs_ready = rhs_load_en;
endmodule
module xls_cmpf32_OGE(
  input wire clk,
  input wire rst,
  input wire [31:0] lhs,
  input wire lhs_valid,
  input wire [31:0] rhs,
  input wire rhs_valid,
  input wire result_ready,
  output wire result,
  output wire result_valid,
  output wire lhs_ready,
  output wire rhs_ready
);
  function automatic priority_sel_1b_3way (input reg [2:0] sel, input reg case0, input reg case1, input reg case2, input reg default_value);
    begin
      casez (sel)
        3'b??1: begin
          priority_sel_1b_3way = case0;
        end
        3'b?10: begin
          priority_sel_1b_3way = case1;
        end
        3'b100: begin
          priority_sel_1b_3way = case2;
        end
        3'b000: begin
          priority_sel_1b_3way = default_value;
        end
        default: begin
          // Propagate X
          priority_sel_1b_3way = 1'dx;
        end
      endcase
    end
  endfunction
  wire [31:0] lhs_reg_init = {1'h0, 8'h00, 23'h00_0000};
  wire [31:0] rhs_reg_init = {1'h0, 8'h00, 23'h00_0000};
  reg [31:0] lhs_reg;
  reg lhs_valid_reg;
  reg [31:0] rhs_reg;
  reg rhs_valid_reg;
  reg result_reg;
  reg result_valid_reg;
  wire [7:0] a_bexp__1;
  wire [7:0] b_bexp__2;
  wire eq_730;
  wire eq_731;
  wire [22:0] a_fraction__2;
  wire [22:0] b_fraction__3;
  wire [22:0] a__1_fraction__5;
  wire [22:0] b__1_fraction__6;
  wire a_sign__2;
  wire b_sign__1;
  wire eq_exp;
  wire gt_fraction;
  wire eq_744;
  wire gt_exp;
  wire and_749;
  wire abs_gt;
  wire result_valid_inv;
  wire p0_all_active_inputs_valid;
  wire result_valid_load_en;
  wire result_load_en;
  wire and_773;
  wire and_774;
  wire p0_stage_done;
  wire lhs_valid_inv;
  wire rhs_valid_inv;
  wire lhs_valid_load_en;
  wire rhs_valid_load_en;
  wire lhs_load_en;
  wire rhs_load_en;
  wire sum;
  assign a_bexp__1 = lhs_reg[30:23];
  assign b_bexp__2 = rhs_reg[30:23];
  assign eq_730 = a_bexp__1 == 8'h00;
  assign eq_731 = b_bexp__2 == 8'h00;
  assign a_fraction__2 = lhs_reg[22:0];
  assign b_fraction__3 = rhs_reg[22:0];
  assign a__1_fraction__5 = a_fraction__2 & {23{~eq_730}};
  assign b__1_fraction__6 = b_fraction__3 & {23{~eq_731}};
  assign a_sign__2 = lhs_reg[31:31];
  assign b_sign__1 = rhs_reg[31:31];
  assign eq_exp = a_bexp__1 == b_bexp__2;
  assign gt_fraction = a__1_fraction__5 > b__1_fraction__6;
  assign eq_744 = a_sign__2 == b_sign__1;
  assign gt_exp = a_bexp__1 > b_bexp__2;
  assign and_749 = eq_730 & eq_731;
  assign abs_gt = gt_exp | eq_exp & gt_fraction;
  assign result_valid_inv = ~result_valid_reg;
  assign p0_all_active_inputs_valid = lhs_valid_reg & rhs_valid_reg;
  assign result_valid_load_en = result_ready | result_valid_inv;
  assign result_load_en = p0_all_active_inputs_valid & result_valid_load_en;
  assign result = priority_sel_1b_3way({~(~a_sign__2 | b_sign__1), ~(a_sign__2 | ~b_sign__1), ~(a_sign__2 | b_sign__1)}, abs_gt, 1'h1, 1'h0, ~abs_gt & ~(eq_744 & eq_exp & a__1_fraction__5 == b__1_fraction__6 | and_749));
  assign and_773 = a_bexp__1 == 8'hff & a_fraction__2 != 23'h00_0000;
  assign and_774 = b_bexp__2 == 8'hff & b_fraction__3 != 23'h00_0000;
  assign p0_stage_done = p0_all_active_inputs_valid & result_load_en;
  assign lhs_valid_inv = ~lhs_valid_reg;
  assign rhs_valid_inv = ~rhs_valid_reg;
  assign lhs_valid_load_en = p0_stage_done | lhs_valid_inv;
  assign rhs_valid_load_en = p0_stage_done | rhs_valid_inv;
  assign lhs_load_en = lhs_valid & lhs_valid_load_en;
  assign rhs_load_en = rhs_valid & rhs_valid_load_en;
  assign sum = ~(and_773 | and_774 | ~result) | ~(and_773 | and_774) & (eq_744 & eq_exp & a_fraction__2 == b_fraction__3 | and_749);
  always @ (posedge clk) begin
    if (rst) begin
      lhs_reg <= lhs_reg_init;
      lhs_valid_reg <= 1'h0;
      rhs_reg <= rhs_reg_init;
      rhs_valid_reg <= 1'h0;
      result_reg <= 1'h0;
      result_valid_reg <= 1'h0;
    end else begin
      lhs_reg <= lhs_load_en ? lhs : lhs_reg;
      lhs_valid_reg <= lhs_valid_load_en ? lhs_valid : lhs_valid_reg;
      rhs_reg <= rhs_load_en ? rhs : rhs_reg;
      rhs_valid_reg <= rhs_valid_load_en ? rhs_valid : rhs_valid_reg;
      result_reg <= result_load_en ? sum : result_reg;
      result_valid_reg <= result_valid_load_en ? p0_all_active_inputs_valid : result_valid_reg;
    end
  end
  assign result = result_reg;
  assign result_valid = result_valid_reg;
  assign lhs_ready = lhs_load_en;
  assign rhs_ready = rhs_load_en;
endmodule
module xls_cmpf32_OGT(
  input wire clk,
  input wire rst,
  input wire [31:0] lhs,
  input wire lhs_valid,
  input wire [31:0] rhs,
  input wire rhs_valid,
  input wire result_ready,
  output wire result,
  output wire result_valid,
  output wire lhs_ready,
  output wire rhs_ready
);
  function automatic priority_sel_1b_3way (input reg [2:0] sel, input reg case0, input reg case1, input reg case2, input reg default_value);
    begin
      casez (sel)
        3'b??1: begin
          priority_sel_1b_3way = case0;
        end
        3'b?10: begin
          priority_sel_1b_3way = case1;
        end
        3'b100: begin
          priority_sel_1b_3way = case2;
        end
        3'b000: begin
          priority_sel_1b_3way = default_value;
        end
        default: begin
          // Propagate X
          priority_sel_1b_3way = 1'dx;
        end
      endcase
    end
  endfunction
  wire [31:0] lhs_reg_init = {1'h0, 8'h00, 23'h00_0000};
  wire [31:0] rhs_reg_init = {1'h0, 8'h00, 23'h00_0000};
  reg [31:0] lhs_reg;
  reg lhs_valid_reg;
  reg [31:0] rhs_reg;
  reg rhs_valid_reg;
  reg result_reg;
  reg result_valid_reg;
  wire [7:0] a_bexp__2;
  wire [7:0] b_bexp__1;
  wire eq_537;
  wire eq_538;
  wire [22:0] a__1_fraction__1;
  wire [22:0] b__1_fraction__2;
  wire eq_exp;
  wire gt_fraction;
  wire a_sign__1;
  wire b_sign;
  wire gt_exp;
  wire result_valid_inv;
  wire abs_gt;
  wire p0_all_active_inputs_valid;
  wire result_valid_load_en;
  wire result_load_en;
  wire p0_stage_done;
  wire lhs_valid_inv;
  wire rhs_valid_inv;
  wire lhs_valid_load_en;
  wire rhs_valid_load_en;
  wire lhs_load_en;
  wire rhs_load_en;
  wire sum;
  assign a_bexp__2 = lhs_reg[30:23];
  assign b_bexp__1 = rhs_reg[30:23];
  assign eq_537 = a_bexp__2 == 8'h00;
  assign eq_538 = b_bexp__1 == 8'h00;
  assign a__1_fraction__1 = lhs_reg[22:0] & {23{~eq_537}};
  assign b__1_fraction__2 = rhs_reg[22:0] & {23{~eq_538}};
  assign eq_exp = a_bexp__2 == b_bexp__1;
  assign gt_fraction = a__1_fraction__1 > b__1_fraction__2;
  assign a_sign__1 = lhs_reg[31:31];
  assign b_sign = rhs_reg[31:31];
  assign gt_exp = a_bexp__2 > b_bexp__1;
  assign result_valid_inv = ~result_valid_reg;
  assign abs_gt = gt_exp | eq_exp & gt_fraction;
  assign p0_all_active_inputs_valid = lhs_valid_reg & rhs_valid_reg;
  assign result_valid_load_en = result_ready | result_valid_inv;
  assign result_load_en = p0_all_active_inputs_valid & result_valid_load_en;
  assign p0_stage_done = p0_all_active_inputs_valid & result_load_en;
  assign lhs_valid_inv = ~lhs_valid_reg;
  assign rhs_valid_inv = ~rhs_valid_reg;
  assign result = priority_sel_1b_3way({~(~a_sign__1 | b_sign), ~(a_sign__1 | ~b_sign), ~(a_sign__1 | b_sign)}, abs_gt, 1'h1, 1'h0, ~abs_gt & ~(eq_exp & a__1_fraction__1 == b__1_fraction__2 | eq_537 & eq_538));
  assign lhs_valid_load_en = p0_stage_done | lhs_valid_inv;
  assign rhs_valid_load_en = p0_stage_done | rhs_valid_inv;
  assign lhs_load_en = lhs_valid & lhs_valid_load_en;
  assign rhs_load_en = rhs_valid & rhs_valid_load_en;
  assign sum = ~(a_bexp__2 == 8'hff & a__1_fraction__1 != 23'h00_0000 | b_bexp__1 == 8'hff & b__1_fraction__2 != 23'h00_0000 | ~result);
  always @ (posedge clk) begin
    if (rst) begin
      lhs_reg <= lhs_reg_init;
      lhs_valid_reg <= 1'h0;
      rhs_reg <= rhs_reg_init;
      rhs_valid_reg <= 1'h0;
      result_reg <= 1'h0;
      result_valid_reg <= 1'h0;
    end else begin
      lhs_reg <= lhs_load_en ? lhs : lhs_reg;
      lhs_valid_reg <= lhs_valid_load_en ? lhs_valid : lhs_valid_reg;
      rhs_reg <= rhs_load_en ? rhs : rhs_reg;
      rhs_valid_reg <= rhs_valid_load_en ? rhs_valid : rhs_valid_reg;
      result_reg <= result_load_en ? sum : result_reg;
      result_valid_reg <= result_valid_load_en ? p0_all_active_inputs_valid : result_valid_reg;
    end
  end
  assign result = result_reg;
  assign result_valid = result_valid_reg;
  assign lhs_ready = lhs_load_en;
  assign rhs_ready = rhs_load_en;
endmodule
module xls_cmpf32_OLE(
  input wire clk,
  input wire rst,
  input wire [31:0] lhs,
  input wire lhs_valid,
  input wire [31:0] rhs,
  input wire rhs_valid,
  input wire result_ready,
  output wire result,
  output wire result_valid,
  output wire lhs_ready,
  output wire rhs_ready
);
  function automatic priority_sel_1b_3way (input reg [2:0] sel, input reg case0, input reg case1, input reg case2, input reg default_value);
    begin
      casez (sel)
        3'b??1: begin
          priority_sel_1b_3way = case0;
        end
        3'b?10: begin
          priority_sel_1b_3way = case1;
        end
        3'b100: begin
          priority_sel_1b_3way = case2;
        end
        3'b000: begin
          priority_sel_1b_3way = default_value;
        end
        default: begin
          // Propagate X
          priority_sel_1b_3way = 1'dx;
        end
      endcase
    end
  endfunction
  wire [31:0] lhs_reg_init = {1'h0, 8'h00, 23'h00_0000};
  wire [31:0] rhs_reg_init = {1'h0, 8'h00, 23'h00_0000};
  reg [31:0] lhs_reg;
  reg lhs_valid_reg;
  reg [31:0] rhs_reg;
  reg rhs_valid_reg;
  reg result_reg;
  reg result_valid_reg;
  wire [7:0] a_bexp__4;
  wire [7:0] b_bexp__2;
  wire eq_695;
  wire eq_696;
  wire [22:0] a_fraction__1;
  wire [22:0] b_fraction;
  wire [22:0] a__1_fraction__5;
  wire [22:0] b__1_fraction__6;
  wire eq_exp;
  wire gt_fraction;
  wire result_valid_inv;
  wire a_sign__2;
  wire b_sign__1;
  wire gt_exp;
  wire p0_all_active_inputs_valid;
  wire result_valid_load_en;
  wire abs_gt;
  wire result_load_en;
  wire p0_stage_done;
  wire lhs_valid_inv;
  wire rhs_valid_inv;
  wire lhs_valid_load_en;
  wire rhs_valid_load_en;
  wire lhs_load_en;
  wire rhs_load_en;
  wire sum;
  assign a_bexp__4 = lhs_reg[30:23];
  assign b_bexp__2 = rhs_reg[30:23];
  assign eq_695 = a_bexp__4 == 8'h00;
  assign eq_696 = b_bexp__2 == 8'h00;
  assign a_fraction__1 = lhs_reg[22:0];
  assign b_fraction = rhs_reg[22:0];
  assign a__1_fraction__5 = a_fraction__1 & {23{~eq_695}};
  assign b__1_fraction__6 = b_fraction & {23{~eq_696}};
  assign eq_exp = a_bexp__4 == b_bexp__2;
  assign gt_fraction = a__1_fraction__5 > b__1_fraction__6;
  assign result_valid_inv = ~result_valid_reg;
  assign a_sign__2 = lhs_reg[31:31];
  assign b_sign__1 = rhs_reg[31:31];
  assign gt_exp = a_bexp__4 > b_bexp__2;
  assign p0_all_active_inputs_valid = lhs_valid_reg & rhs_valid_reg;
  assign result_valid_load_en = result_ready | result_valid_inv;
  assign abs_gt = gt_exp | eq_exp & gt_fraction;
  assign result_load_en = p0_all_active_inputs_valid & result_valid_load_en;
  assign p0_stage_done = p0_all_active_inputs_valid & result_load_en;
  assign lhs_valid_inv = ~lhs_valid_reg;
  assign rhs_valid_inv = ~rhs_valid_reg;
  assign lhs_valid_load_en = p0_stage_done | lhs_valid_inv;
  assign rhs_valid_load_en = p0_stage_done | rhs_valid_inv;
  assign result = priority_sel_1b_3way({~(~a_sign__2 | b_sign__1), ~(a_sign__2 | ~b_sign__1), ~(a_sign__2 | b_sign__1)}, abs_gt, 1'h1, 1'h0, ~abs_gt & ~(eq_exp & a__1_fraction__5 == b__1_fraction__6 | eq_695 & eq_696));
  assign lhs_load_en = lhs_valid & lhs_valid_load_en;
  assign rhs_load_en = rhs_valid & rhs_valid_load_en;
  assign sum = ~(a_bexp__4 == 8'hff & a_fraction__1 != 23'h00_0000 | b_bexp__2 == 8'hff & b_fraction != 23'h00_0000 | result);
  always @ (posedge clk) begin
    if (rst) begin
      lhs_reg <= lhs_reg_init;
      lhs_valid_reg <= 1'h0;
      rhs_reg <= rhs_reg_init;
      rhs_valid_reg <= 1'h0;
      result_reg <= 1'h0;
      result_valid_reg <= 1'h0;
    end else begin
      lhs_reg <= lhs_load_en ? lhs : lhs_reg;
      lhs_valid_reg <= lhs_valid_load_en ? lhs_valid : lhs_valid_reg;
      rhs_reg <= rhs_load_en ? rhs : rhs_reg;
      rhs_valid_reg <= rhs_valid_load_en ? rhs_valid : rhs_valid_reg;
      result_reg <= result_load_en ? sum : result_reg;
      result_valid_reg <= result_valid_load_en ? p0_all_active_inputs_valid : result_valid_reg;
    end
  end
  assign result = result_reg;
  assign result_valid = result_valid_reg;
  assign lhs_ready = lhs_load_en;
  assign rhs_ready = rhs_load_en;
endmodule
module xls_cmpf32_OLT(
  input wire clk,
  input wire rst,
  input wire [31:0] lhs,
  input wire lhs_valid,
  input wire [31:0] rhs,
  input wire rhs_valid,
  input wire result_ready,
  output wire result,
  output wire result_valid,
  output wire lhs_ready,
  output wire rhs_ready
);
  function automatic priority_sel_1b_3way (input reg [2:0] sel, input reg case0, input reg case1, input reg case2, input reg default_value);
    begin
      casez (sel)
        3'b??1: begin
          priority_sel_1b_3way = case0;
        end
        3'b?10: begin
          priority_sel_1b_3way = case1;
        end
        3'b100: begin
          priority_sel_1b_3way = case2;
        end
        3'b000: begin
          priority_sel_1b_3way = default_value;
        end
        default: begin
          // Propagate X
          priority_sel_1b_3way = 1'dx;
        end
      endcase
    end
  endfunction
  wire [31:0] lhs_reg_init = {1'h0, 8'h00, 23'h00_0000};
  wire [31:0] rhs_reg_init = {1'h0, 8'h00, 23'h00_0000};
  reg [31:0] lhs_reg;
  reg lhs_valid_reg;
  reg [31:0] rhs_reg;
  reg rhs_valid_reg;
  reg result_reg;
  reg result_valid_reg;
  wire [7:0] a_bexp__4;
  wire [7:0] b_bexp__1;
  wire eq_923;
  wire eq_924;
  wire [22:0] a_fraction__5;
  wire [22:0] b_fraction__4;
  wire [22:0] a__1_fraction__1;
  wire [22:0] b__1_fraction__2;
  wire eq_exp;
  wire gt_fraction;
  wire a_sign__1;
  wire b_sign__2;
  wire gt_exp;
  wire result_valid_inv;
  wire abs_gt;
  wire eq_942;
  wire p0_all_active_inputs_valid;
  wire result_valid_load_en;
  wire result_load_en;
  wire p0_stage_done;
  wire lhs_valid_inv;
  wire rhs_valid_inv;
  wire lhs_valid_load_en;
  wire rhs_valid_load_en;
  wire lhs_load_en;
  wire rhs_load_en;
  wire sum;
  assign a_bexp__4 = lhs_reg[30:23];
  assign b_bexp__1 = rhs_reg[30:23];
  assign eq_923 = a_bexp__4 == 8'h00;
  assign eq_924 = b_bexp__1 == 8'h00;
  assign a_fraction__5 = lhs_reg[22:0];
  assign b_fraction__4 = rhs_reg[22:0];
  assign a__1_fraction__1 = a_fraction__5 & {23{~eq_923}};
  assign b__1_fraction__2 = b_fraction__4 & {23{~eq_924}};
  assign eq_exp = a_bexp__4 == b_bexp__1;
  assign gt_fraction = a__1_fraction__1 > b__1_fraction__2;
  assign a_sign__1 = lhs_reg[31:31];
  assign b_sign__2 = rhs_reg[31:31];
  assign gt_exp = a_bexp__4 > b_bexp__1;
  assign result_valid_inv = ~result_valid_reg;
  assign abs_gt = gt_exp | eq_exp & gt_fraction;
  assign eq_942 = a_sign__1 == b_sign__2;
  assign p0_all_active_inputs_valid = lhs_valid_reg & rhs_valid_reg;
  assign result_valid_load_en = result_ready | result_valid_inv;
  assign result_load_en = p0_all_active_inputs_valid & result_valid_load_en;
  assign p0_stage_done = p0_all_active_inputs_valid & result_load_en;
  assign lhs_valid_inv = ~lhs_valid_reg;
  assign rhs_valid_inv = ~rhs_valid_reg;
  assign result = priority_sel_1b_3way({~(~a_sign__1 | b_sign__2), ~(a_sign__1 | ~b_sign__2), ~(a_sign__1 | b_sign__2)}, abs_gt, 1'h1, 1'h0, ~abs_gt & ~(eq_942 & eq_exp & a__1_fraction__1 == b__1_fraction__2));
  assign lhs_valid_load_en = p0_stage_done | lhs_valid_inv;
  assign rhs_valid_load_en = p0_stage_done | rhs_valid_inv;
  assign lhs_load_en = lhs_valid & lhs_valid_load_en;
  assign rhs_load_en = rhs_valid & rhs_valid_load_en;
  assign sum = ~(a_bexp__4 == 8'hff & a_fraction__5 != 23'h00_0000 | b_bexp__1 == 8'hff & b_fraction__4 != 23'h00_0000 | (result | eq_942 & eq_exp & a_fraction__5 == b_fraction__4 | eq_923 & eq_924));
  always @ (posedge clk) begin
    if (rst) begin
      lhs_reg <= lhs_reg_init;
      lhs_valid_reg <= 1'h0;
      rhs_reg <= rhs_reg_init;
      rhs_valid_reg <= 1'h0;
      result_reg <= 1'h0;
      result_valid_reg <= 1'h0;
    end else begin
      lhs_reg <= lhs_load_en ? lhs : lhs_reg;
      lhs_valid_reg <= lhs_valid_load_en ? lhs_valid : lhs_valid_reg;
      rhs_reg <= rhs_load_en ? rhs : rhs_reg;
      rhs_valid_reg <= rhs_valid_load_en ? rhs_valid : rhs_valid_reg;
      result_reg <= result_load_en ? sum : result_reg;
      result_valid_reg <= result_valid_load_en ? p0_all_active_inputs_valid : result_valid_reg;
    end
  end
  assign result = result_reg;
  assign result_valid = result_valid_reg;
  assign lhs_ready = lhs_load_en;
  assign rhs_ready = rhs_load_en;
endmodule
module xls_divf32(
  input wire clk,
  input wire rst,
  input wire [31:0] lhs,
  input wire lhs_valid,
  input wire [31:0] rhs,
  input wire rhs_valid,
  input wire result_ready,
  output wire [31:0] result,
  output wire result_valid,
  output wire lhs_ready,
  output wire rhs_ready
);
  wire [31:0] lhs_reg_init = {1'h0, 8'h00, 23'h00_0000};
  wire [31:0] rhs_reg_init = {1'h0, 8'h00, 23'h00_0000};
  wire [31:0] result_reg_init = {1'h0, 8'h00, 23'h00_0000};
  reg p0_bit_slice_3967;
  reg p0_bit_slice_3968;
  reg p0_bit_slice_3969;
  reg p0_bit_slice_3970;
  reg p0_bit_slice_3971;
  reg p0_bit_slice_3972;
  reg p0_bit_slice_3973;
  reg p0_bit_slice_3974;
  reg p0_bit_slice_3975;
  reg p0_bit_slice_3976;
  reg p0_bit_slice_3977;
  reg p0_bit_slice_3978;
  reg p0_bit_slice_3979;
  reg p0_bit_slice_3980;
  reg p0_bit_slice_3981;
  reg p0_bit_slice_3982;
  reg p0_bit_slice_3983;
  reg p0_bit_slice_3984;
  reg p0_bit_slice_3985;
  reg p0_bit_slice_3986;
  reg p0_bit_slice_3987;
  reg [7:0] p0_a_bexp;
  reg p0_bit_slice_3989;
  reg p0_bit_slice_3990;
  reg p0_a_sign;
  reg [22:0] p1_concat_4053;
  reg [22:0] p1_b_fraction;
  reg p1_bit_slice_3968;
  reg p1_bit_slice_3969;
  reg p1_bit_slice_3970;
  reg p1_bit_slice_3971;
  reg p1_bit_slice_3972;
  reg p1_bit_slice_3973;
  reg p1_bit_slice_3974;
  reg p1_bit_slice_3975;
  reg p1_bit_slice_3976;
  reg p1_bit_slice_3977;
  reg p1_bit_slice_3978;
  reg p1_bit_slice_3979;
  reg p1_bit_slice_3980;
  reg p1_bit_slice_3981;
  reg p1_bit_slice_3982;
  reg p1_bit_slice_3983;
  reg p1_bit_slice_3984;
  reg p1_bit_slice_3985;
  reg p1_bit_slice_3986;
  reg p1_bit_slice_3987;
  reg [7:0] p1_a_bexp;
  reg [7:0] p1_b_bexp;
  reg p1_bit_slice_3989;
  reg p1_bit_slice_3990;
  reg p1_result_sign;
  reg [22:0] p2_b_fraction;
  reg p2_uge_4116;
  reg [23:0] p2_b_fractionivisor__1;
  reg [22:0] p2_concat_4123;
  reg p2_uge_4124;
  reg p2_bit_slice_3969;
  reg p2_bit_slice_3970;
  reg p2_bit_slice_3971;
  reg p2_bit_slice_3972;
  reg p2_bit_slice_3973;
  reg p2_bit_slice_3974;
  reg p2_bit_slice_3975;
  reg p2_bit_slice_3976;
  reg p2_bit_slice_3977;
  reg p2_bit_slice_3978;
  reg p2_bit_slice_3979;
  reg p2_bit_slice_3980;
  reg p2_bit_slice_3981;
  reg p2_bit_slice_3982;
  reg p2_bit_slice_3983;
  reg p2_bit_slice_3984;
  reg p2_bit_slice_3985;
  reg p2_bit_slice_3986;
  reg p2_bit_slice_3987;
  reg p2_bit_slice_3989;
  reg [8:0] p2_signed_exp_s9;
  reg p2_bit_slice_3990;
  reg p2_result_sign;
  reg [22:0] p3_b_fraction;
  reg p3_uge_4116;
  reg [23:0] p3_b_fractionivisor__1;
  reg p3_uge_4124;
  reg [22:0] p3_concat_4194;
  reg p3_uge_4195;
  reg p3_bit_slice_3970;
  reg p3_bit_slice_3971;
  reg p3_bit_slice_3972;
  reg p3_bit_slice_3973;
  reg p3_bit_slice_3974;
  reg p3_bit_slice_3975;
  reg p3_bit_slice_3976;
  reg p3_bit_slice_3977;
  reg p3_bit_slice_3978;
  reg p3_bit_slice_3979;
  reg p3_bit_slice_3980;
  reg p3_bit_slice_3981;
  reg p3_bit_slice_3982;
  reg p3_bit_slice_3983;
  reg p3_bit_slice_3984;
  reg p3_bit_slice_3985;
  reg p3_bit_slice_3986;
  reg p3_bit_slice_3987;
  reg p3_bit_slice_3989;
  reg p3_bit_slice_3990;
  reg p3_flag_zero;
  reg p3_result_sign;
  reg [7:0] p3_result_exp;
  reg [22:0] p4_b_fraction;
  reg p4_uge_4116;
  reg [23:0] p4_b_fractionivisor__1;
  reg p4_uge_4124;
  reg p4_uge_4195;
  reg [22:0] p4_concat_4269;
  reg p4_uge_4270;
  reg p4_bit_slice_3971;
  reg p4_bit_slice_3972;
  reg p4_bit_slice_3973;
  reg p4_bit_slice_3974;
  reg p4_bit_slice_3975;
  reg p4_bit_slice_3976;
  reg p4_bit_slice_3977;
  reg p4_bit_slice_3978;
  reg p4_bit_slice_3979;
  reg p4_bit_slice_3980;
  reg p4_bit_slice_3981;
  reg p4_bit_slice_3982;
  reg p4_bit_slice_3983;
  reg p4_bit_slice_3984;
  reg p4_bit_slice_3985;
  reg p4_bit_slice_3986;
  reg p4_bit_slice_3987;
  reg p4_bit_slice_3989;
  reg p4_bit_slice_3990;
  reg p4_flag_zero;
  reg p4_result_sign;
  reg [7:0] p4_result_exp;
  reg [22:0] p5_b_fraction;
  reg p5_uge_4116;
  reg [23:0] p5_b_fractionivisor__1;
  reg p5_uge_4124;
  reg p5_uge_4195;
  reg p5_uge_4270;
  reg [22:0] p5_concat_4335;
  reg p5_uge_4336;
  reg p5_bit_slice_3972;
  reg p5_bit_slice_3973;
  reg p5_bit_slice_3974;
  reg p5_bit_slice_3975;
  reg p5_bit_slice_3976;
  reg p5_bit_slice_3977;
  reg p5_bit_slice_3978;
  reg p5_bit_slice_3979;
  reg p5_bit_slice_3980;
  reg p5_bit_slice_3981;
  reg p5_bit_slice_3982;
  reg p5_bit_slice_3983;
  reg p5_bit_slice_3984;
  reg p5_bit_slice_3985;
  reg p5_bit_slice_3986;
  reg p5_bit_slice_3987;
  reg p5_bit_slice_3989;
  reg p5_bit_slice_3990;
  reg p5_flag_zero;
  reg p5_result_sign;
  reg [7:0] p5_result_exp;
  reg [22:0] p6_b_fraction;
  reg p6_uge_4116;
  reg [23:0] p6_b_fractionivisor__1;
  reg p6_uge_4124;
  reg p6_uge_4195;
  reg p6_uge_4270;
  reg p6_uge_4336;
  reg [22:0] p6_concat_4401;
  reg p6_uge_4402;
  reg p6_bit_slice_3973;
  reg p6_bit_slice_3974;
  reg p6_bit_slice_3975;
  reg p6_bit_slice_3976;
  reg p6_bit_slice_3977;
  reg p6_bit_slice_3978;
  reg p6_bit_slice_3979;
  reg p6_bit_slice_3980;
  reg p6_bit_slice_3981;
  reg p6_bit_slice_3982;
  reg p6_bit_slice_3983;
  reg p6_bit_slice_3984;
  reg p6_bit_slice_3985;
  reg p6_bit_slice_3986;
  reg p6_bit_slice_3987;
  reg p6_bit_slice_3989;
  reg p6_bit_slice_3990;
  reg p6_flag_zero;
  reg p6_result_sign;
  reg [7:0] p6_result_exp;
  reg [22:0] p7_b_fraction;
  reg p7_uge_4116;
  reg [23:0] p7_b_fractionivisor__1;
  reg p7_uge_4124;
  reg p7_uge_4195;
  reg p7_uge_4270;
  reg p7_uge_4336;
  reg p7_uge_4402;
  reg [22:0] p7_concat_4467;
  reg p7_uge_4468;
  reg p7_bit_slice_3974;
  reg p7_bit_slice_3975;
  reg p7_bit_slice_3976;
  reg p7_bit_slice_3977;
  reg p7_bit_slice_3978;
  reg p7_bit_slice_3979;
  reg p7_bit_slice_3980;
  reg p7_bit_slice_3981;
  reg p7_bit_slice_3982;
  reg p7_bit_slice_3983;
  reg p7_bit_slice_3984;
  reg p7_bit_slice_3985;
  reg p7_bit_slice_3986;
  reg p7_bit_slice_3987;
  reg p7_bit_slice_3989;
  reg p7_bit_slice_3990;
  reg p7_flag_zero;
  reg p7_result_sign;
  reg [7:0] p7_result_exp;
  reg [22:0] p8_b_fraction;
  reg p8_uge_4116;
  reg [23:0] p8_b_fractionivisor__1;
  reg p8_uge_4124;
  reg p8_uge_4195;
  reg p8_uge_4270;
  reg p8_uge_4336;
  reg p8_uge_4402;
  reg p8_uge_4468;
  reg [22:0] p8_concat_4533;
  reg p8_uge_4534;
  reg p8_bit_slice_3975;
  reg p8_bit_slice_3976;
  reg p8_bit_slice_3977;
  reg p8_bit_slice_3978;
  reg p8_bit_slice_3979;
  reg p8_bit_slice_3980;
  reg p8_bit_slice_3981;
  reg p8_bit_slice_3982;
  reg p8_bit_slice_3983;
  reg p8_bit_slice_3984;
  reg p8_bit_slice_3985;
  reg p8_bit_slice_3986;
  reg p8_bit_slice_3987;
  reg p8_bit_slice_3989;
  reg p8_bit_slice_3990;
  reg p8_flag_zero;
  reg p8_result_sign;
  reg [7:0] p8_result_exp;
  reg [22:0] p9_b_fraction;
  reg p9_uge_4116;
  reg [23:0] p9_b_fractionivisor__1;
  reg p9_uge_4124;
  reg p9_uge_4195;
  reg p9_uge_4270;
  reg p9_uge_4336;
  reg p9_uge_4402;
  reg p9_uge_4468;
  reg p9_uge_4534;
  reg [22:0] p9_concat_4599;
  reg p9_uge_4600;
  reg p9_bit_slice_3976;
  reg p9_bit_slice_3977;
  reg p9_bit_slice_3978;
  reg p9_bit_slice_3979;
  reg p9_bit_slice_3980;
  reg p9_bit_slice_3981;
  reg p9_bit_slice_3982;
  reg p9_bit_slice_3983;
  reg p9_bit_slice_3984;
  reg p9_bit_slice_3985;
  reg p9_bit_slice_3986;
  reg p9_bit_slice_3987;
  reg p9_bit_slice_3989;
  reg p9_bit_slice_3990;
  reg p9_flag_zero;
  reg p9_result_sign;
  reg [7:0] p9_result_exp;
  reg [22:0] p10_b_fraction;
  reg p10_uge_4116;
  reg [23:0] p10_b_fractionivisor__1;
  reg p10_uge_4124;
  reg p10_uge_4195;
  reg p10_uge_4270;
  reg p10_uge_4336;
  reg p10_uge_4402;
  reg p10_uge_4468;
  reg p10_uge_4534;
  reg p10_uge_4600;
  reg [22:0] p10_concat_4665;
  reg p10_uge_4666;
  reg p10_bit_slice_3977;
  reg p10_bit_slice_3978;
  reg p10_bit_slice_3979;
  reg p10_bit_slice_3980;
  reg p10_bit_slice_3981;
  reg p10_bit_slice_3982;
  reg p10_bit_slice_3983;
  reg p10_bit_slice_3984;
  reg p10_bit_slice_3985;
  reg p10_bit_slice_3986;
  reg p10_bit_slice_3987;
  reg p10_bit_slice_3989;
  reg p10_bit_slice_3990;
  reg p10_flag_zero;
  reg p10_result_sign;
  reg [7:0] p10_result_exp;
  reg [22:0] p11_b_fraction;
  reg p11_uge_4116;
  reg [23:0] p11_b_fractionivisor__1;
  reg p11_uge_4124;
  reg p11_uge_4195;
  reg p11_uge_4270;
  reg p11_uge_4336;
  reg p11_uge_4402;
  reg p11_uge_4468;
  reg p11_uge_4534;
  reg p11_uge_4600;
  reg p11_uge_4666;
  reg [22:0] p11_concat_4731;
  reg p11_uge_4732;
  reg p11_bit_slice_3978;
  reg p11_bit_slice_3979;
  reg p11_bit_slice_3980;
  reg p11_bit_slice_3981;
  reg p11_bit_slice_3982;
  reg p11_bit_slice_3983;
  reg p11_bit_slice_3984;
  reg p11_bit_slice_3985;
  reg p11_bit_slice_3986;
  reg p11_bit_slice_3987;
  reg p11_bit_slice_3989;
  reg p11_bit_slice_3990;
  reg p11_flag_zero;
  reg p11_result_sign;
  reg [7:0] p11_result_exp;
  reg [22:0] p12_b_fraction;
  reg p12_uge_4116;
  reg [23:0] p12_b_fractionivisor__1;
  reg p12_uge_4124;
  reg p12_uge_4195;
  reg p12_uge_4270;
  reg p12_uge_4336;
  reg p12_uge_4402;
  reg p12_uge_4468;
  reg p12_uge_4534;
  reg p12_uge_4600;
  reg p12_uge_4666;
  reg p12_uge_4732;
  reg [22:0] p12_concat_4797;
  reg p12_uge_4798;
  reg p12_bit_slice_3979;
  reg p12_bit_slice_3980;
  reg p12_bit_slice_3981;
  reg p12_bit_slice_3982;
  reg p12_bit_slice_3983;
  reg p12_bit_slice_3984;
  reg p12_bit_slice_3985;
  reg p12_bit_slice_3986;
  reg p12_bit_slice_3987;
  reg p12_bit_slice_3989;
  reg p12_bit_slice_3990;
  reg p12_flag_zero;
  reg p12_result_sign;
  reg [7:0] p12_result_exp;
  reg [22:0] p13_b_fraction;
  reg p13_uge_4116;
  reg [23:0] p13_b_fractionivisor__1;
  reg p13_uge_4124;
  reg p13_uge_4195;
  reg p13_uge_4270;
  reg p13_uge_4336;
  reg p13_uge_4402;
  reg p13_uge_4468;
  reg p13_uge_4534;
  reg p13_uge_4600;
  reg p13_uge_4666;
  reg p13_uge_4732;
  reg p13_uge_4798;
  reg [22:0] p13_concat_4863;
  reg p13_uge_4864;
  reg p13_bit_slice_3980;
  reg p13_bit_slice_3981;
  reg p13_bit_slice_3982;
  reg p13_bit_slice_3983;
  reg p13_bit_slice_3984;
  reg p13_bit_slice_3985;
  reg p13_bit_slice_3986;
  reg p13_bit_slice_3987;
  reg p13_bit_slice_3989;
  reg p13_bit_slice_3990;
  reg p13_flag_zero;
  reg p13_result_sign;
  reg [7:0] p13_result_exp;
  reg [22:0] p14_b_fraction;
  reg p14_uge_4116;
  reg [23:0] p14_b_fractionivisor__1;
  reg p14_uge_4124;
  reg p14_uge_4195;
  reg p14_uge_4270;
  reg p14_uge_4336;
  reg p14_uge_4402;
  reg p14_uge_4468;
  reg p14_uge_4534;
  reg p14_uge_4600;
  reg p14_uge_4666;
  reg p14_uge_4732;
  reg p14_uge_4798;
  reg p14_uge_4864;
  reg [22:0] p14_concat_4929;
  reg p14_uge_4930;
  reg p14_bit_slice_3981;
  reg p14_bit_slice_3982;
  reg p14_bit_slice_3983;
  reg p14_bit_slice_3984;
  reg p14_bit_slice_3985;
  reg p14_bit_slice_3986;
  reg p14_bit_slice_3987;
  reg p14_bit_slice_3989;
  reg p14_bit_slice_3990;
  reg p14_flag_zero;
  reg p14_result_sign;
  reg [7:0] p14_result_exp;
  reg [22:0] p15_b_fraction;
  reg p15_uge_4116;
  reg [23:0] p15_b_fractionivisor__1;
  reg p15_uge_4124;
  reg p15_uge_4195;
  reg p15_uge_4270;
  reg p15_uge_4336;
  reg p15_uge_4402;
  reg p15_uge_4468;
  reg p15_uge_4534;
  reg p15_uge_4600;
  reg p15_uge_4666;
  reg p15_uge_4732;
  reg p15_uge_4798;
  reg p15_uge_4864;
  reg p15_uge_4930;
  reg [22:0] p15_concat_4995;
  reg p15_uge_4996;
  reg p15_bit_slice_3982;
  reg p15_bit_slice_3983;
  reg p15_bit_slice_3984;
  reg p15_bit_slice_3985;
  reg p15_bit_slice_3986;
  reg p15_bit_slice_3987;
  reg p15_bit_slice_3989;
  reg p15_bit_slice_3990;
  reg p15_flag_zero;
  reg p15_result_sign;
  reg [7:0] p15_result_exp;
  reg [22:0] p16_b_fraction;
  reg p16_uge_4116;
  reg [23:0] p16_b_fractionivisor__1;
  reg p16_uge_4124;
  reg p16_uge_4195;
  reg p16_uge_4270;
  reg p16_uge_4336;
  reg p16_uge_4402;
  reg p16_uge_4468;
  reg p16_uge_4534;
  reg p16_uge_4600;
  reg p16_uge_4666;
  reg p16_uge_4732;
  reg p16_uge_4798;
  reg p16_uge_4864;
  reg p16_uge_4930;
  reg p16_uge_4996;
  reg [22:0] p16_concat_5061;
  reg p16_uge_5062;
  reg p16_bit_slice_3983;
  reg p16_bit_slice_3984;
  reg p16_bit_slice_3985;
  reg p16_bit_slice_3986;
  reg p16_bit_slice_3987;
  reg p16_bit_slice_3989;
  reg p16_bit_slice_3990;
  reg p16_flag_zero;
  reg p16_result_sign;
  reg [7:0] p16_result_exp;
  reg [22:0] p17_b_fraction;
  reg p17_uge_4116;
  reg [23:0] p17_b_fractionivisor__1;
  reg p17_uge_4124;
  reg p17_uge_4195;
  reg p17_uge_4270;
  reg p17_uge_4336;
  reg p17_uge_4402;
  reg p17_uge_4468;
  reg p17_uge_4534;
  reg p17_uge_4600;
  reg p17_uge_4666;
  reg p17_uge_4732;
  reg p17_uge_4798;
  reg p17_uge_4864;
  reg p17_uge_4930;
  reg p17_uge_4996;
  reg p17_uge_5062;
  reg [22:0] p17_concat_5127;
  reg p17_uge_5128;
  reg p17_bit_slice_3984;
  reg p17_bit_slice_3985;
  reg p17_bit_slice_3986;
  reg p17_bit_slice_3987;
  reg p17_bit_slice_3989;
  reg p17_bit_slice_3990;
  reg p17_flag_zero;
  reg p17_result_sign;
  reg [7:0] p17_result_exp;
  reg [22:0] p18_b_fraction;
  reg p18_uge_4116;
  reg [23:0] p18_b_fractionivisor__1;
  reg p18_uge_4124;
  reg p18_uge_4195;
  reg p18_uge_4270;
  reg p18_uge_4336;
  reg p18_uge_4402;
  reg p18_uge_4468;
  reg p18_uge_4534;
  reg p18_uge_4600;
  reg p18_uge_4666;
  reg p18_uge_4732;
  reg p18_uge_4798;
  reg p18_uge_4864;
  reg p18_uge_4930;
  reg p18_uge_4996;
  reg p18_uge_5062;
  reg p18_uge_5128;
  reg [22:0] p18_concat_5193;
  reg p18_uge_5194;
  reg p18_bit_slice_3985;
  reg p18_bit_slice_3986;
  reg p18_bit_slice_3987;
  reg p18_bit_slice_3989;
  reg p18_bit_slice_3990;
  reg p18_flag_zero;
  reg p18_result_sign;
  reg [7:0] p18_result_exp;
  reg [22:0] p19_b_fraction;
  reg p19_uge_4116;
  reg [23:0] p19_b_fractionivisor__1;
  reg p19_uge_4124;
  reg p19_uge_4195;
  reg p19_uge_4270;
  reg p19_uge_4336;
  reg p19_uge_4402;
  reg p19_uge_4468;
  reg p19_uge_4534;
  reg p19_uge_4600;
  reg p19_uge_4666;
  reg p19_uge_4732;
  reg p19_uge_4798;
  reg p19_uge_4864;
  reg p19_uge_4930;
  reg p19_uge_4996;
  reg p19_uge_5062;
  reg p19_uge_5128;
  reg p19_uge_5194;
  reg [22:0] p19_concat_5259;
  reg p19_uge_5260;
  reg p19_bit_slice_3986;
  reg p19_bit_slice_3987;
  reg p19_bit_slice_3989;
  reg p19_bit_slice_3990;
  reg p19_flag_zero;
  reg p19_result_sign;
  reg [7:0] p19_result_exp;
  reg [22:0] p20_b_fraction;
  reg p20_uge_4116;
  reg [23:0] p20_b_fractionivisor__1;
  reg p20_uge_4124;
  reg p20_uge_4195;
  reg p20_uge_4270;
  reg p20_uge_4336;
  reg p20_uge_4402;
  reg p20_uge_4468;
  reg p20_uge_4534;
  reg p20_uge_4600;
  reg p20_uge_4666;
  reg p20_uge_4732;
  reg p20_uge_4798;
  reg p20_uge_4864;
  reg p20_uge_4930;
  reg p20_uge_4996;
  reg p20_uge_5062;
  reg p20_uge_5128;
  reg p20_uge_5194;
  reg p20_uge_5260;
  reg [22:0] p20_concat_5325;
  reg p20_uge_5326;
  reg p20_bit_slice_3987;
  reg p20_bit_slice_3989;
  reg p20_bit_slice_3990;
  reg p20_flag_zero;
  reg p20_result_sign;
  reg [7:0] p20_result_exp;
  reg [22:0] p21_b_fraction;
  reg p21_uge_4116;
  reg [23:0] p21_b_fractionivisor__1;
  reg p21_uge_4124;
  reg p21_uge_4195;
  reg p21_uge_4270;
  reg p21_uge_4336;
  reg p21_uge_4402;
  reg p21_uge_4468;
  reg p21_uge_4534;
  reg p21_uge_4600;
  reg p21_uge_4666;
  reg p21_uge_4732;
  reg p21_uge_4798;
  reg p21_uge_4864;
  reg p21_uge_4930;
  reg p21_uge_4996;
  reg p21_uge_5062;
  reg p21_uge_5128;
  reg p21_uge_5194;
  reg p21_uge_5260;
  reg p21_uge_5326;
  reg [22:0] p21_concat_5391;
  reg p21_uge_5392;
  reg p21_bit_slice_3989;
  reg p21_bit_slice_3990;
  reg p21_flag_zero;
  reg p21_result_sign;
  reg [7:0] p21_result_exp;
  reg [22:0] p22_b_fraction;
  reg p22_uge_4116;
  reg [23:0] p22_b_fractionivisor__1;
  reg p22_uge_4124;
  reg p22_uge_4195;
  reg p22_uge_4270;
  reg p22_uge_4336;
  reg p22_uge_4402;
  reg p22_uge_4468;
  reg p22_uge_4534;
  reg p22_uge_4600;
  reg p22_uge_4666;
  reg p22_uge_4732;
  reg p22_uge_4798;
  reg p22_uge_4864;
  reg p22_uge_4930;
  reg p22_uge_4996;
  reg p22_uge_5062;
  reg p22_uge_5128;
  reg p22_uge_5194;
  reg p22_uge_5260;
  reg p22_uge_5326;
  reg p22_uge_5392;
  reg [22:0] p22_concat_5457;
  reg p22_uge_5458;
  reg p22_bit_slice_3990;
  reg p22_flag_zero;
  reg p22_result_sign;
  reg [7:0] p22_result_exp;
  reg p23_uge_4116;
  reg p23_uge_4124;
  reg p23_uge_4195;
  reg p23_uge_4270;
  reg p23_uge_4336;
  reg p23_uge_4402;
  reg p23_uge_4468;
  reg p23_uge_4534;
  reg p23_uge_4600;
  reg p23_uge_4666;
  reg p23_uge_4732;
  reg p23_uge_4798;
  reg p23_uge_4864;
  reg p23_uge_4930;
  reg p23_uge_4996;
  reg p23_uge_5062;
  reg p23_uge_5128;
  reg p23_uge_5194;
  reg p23_uge_5260;
  reg p23_uge_5326;
  reg p23_uge_5392;
  reg p23_uge_5458;
  reg p23_flag_zero;
  reg p23_q__23_squeezed_portion_0_width_1;
  reg p23_result_sign;
  reg [7:0] p23_result_exp;
  reg p0_valid;
  reg p1_valid;
  reg p2_valid;
  reg p3_valid;
  reg p4_valid;
  reg p5_valid;
  reg p6_valid;
  reg p7_valid;
  reg p8_valid;
  reg p9_valid;
  reg p10_valid;
  reg p11_valid;
  reg p12_valid;
  reg p13_valid;
  reg p14_valid;
  reg p15_valid;
  reg p16_valid;
  reg p17_valid;
  reg p18_valid;
  reg p19_valid;
  reg p20_valid;
  reg p21_valid;
  reg p22_valid;
  reg p23_valid;
  reg p24_valid;
  reg p25_valid;
  reg p26_valid;
  reg p27_valid;
  reg p28_valid;
  reg p29_valid;
  reg p30_valid;
  reg [31:0] lhs_reg;
  reg lhs_valid_reg;
  reg [31:0] rhs_reg;
  reg rhs_valid_reg;
  reg [31:0] result_reg;
  reg result_valid_reg;
  wire result_valid_inv;
  wire result_valid_load_en;
  wire result_load_en;
  wire p24_stage_done;
  wire p24_not_valid;
  wire p23_enable;
  wire p23_data_enable;
  wire p23_not_valid;
  wire p22_enable;
  wire p22_data_enable;
  wire p22_not_valid;
  wire p21_enable;
  wire p21_data_enable;
  wire p21_not_valid;
  wire p20_enable;
  wire p20_data_enable;
  wire p20_not_valid;
  wire p19_enable;
  wire p19_data_enable;
  wire p19_not_valid;
  wire p18_enable;
  wire p18_data_enable;
  wire p18_not_valid;
  wire p17_enable;
  wire p17_data_enable;
  wire p17_not_valid;
  wire p16_enable;
  wire p16_data_enable;
  wire p16_not_valid;
  wire p15_enable;
  wire p15_data_enable;
  wire p15_not_valid;
  wire p14_enable;
  wire p14_data_enable;
  wire p14_not_valid;
  wire p13_enable;
  wire p13_data_enable;
  wire p13_not_valid;
  wire p12_enable;
  wire p12_data_enable;
  wire p12_not_valid;
  wire p11_enable;
  wire p11_data_enable;
  wire p11_not_valid;
  wire p10_enable;
  wire p10_data_enable;
  wire p10_not_valid;
  wire p9_enable;
  wire p9_data_enable;
  wire p9_not_valid;
  wire p8_enable;
  wire p8_data_enable;
  wire p8_not_valid;
  wire p7_enable;
  wire p7_data_enable;
  wire p7_not_valid;
  wire p6_enable;
  wire p6_data_enable;
  wire p6_not_valid;
  wire p5_enable;
  wire p5_data_enable;
  wire p5_not_valid;
  wire p4_enable;
  wire p4_data_enable;
  wire p4_not_valid;
  wire p3_enable;
  wire p3_data_enable;
  wire p3_not_valid;
  wire p2_enable;
  wire p2_data_enable;
  wire p2_not_valid;
  wire p1_enable;
  wire p1_stage_done;
  wire p1_data_enable;
  wire p1_not_valid;
  wire [22:0] sub_5519;
  wire [22:0] sub_5453;
  wire [22:0] sub_5387;
  wire [22:0] sub_5321;
  wire [22:0] sub_5255;
  wire [22:0] sub_5189;
  wire [22:0] sub_5123;
  wire [22:0] sub_5057;
  wire [22:0] sub_4991;
  wire [22:0] sub_4925;
  wire [22:0] sub_4859;
  wire [22:0] sub_4793;
  wire [22:0] sub_4727;
  wire [22:0] sub_4661;
  wire [22:0] sub_4595;
  wire [22:0] sub_4529;
  wire [22:0] sub_4463;
  wire [22:0] sub_4397;
  wire [22:0] sub_4331;
  wire [22:0] sub_4265;
  wire [22:0] sub_4190;
  wire flag_zero;
  wire uge_4116;
  wire [22:0] sub_4117;
  wire p0_enable;
  wire [22:0] r__68;
  wire [22:0] r__67;
  wire [22:0] r__66;
  wire [22:0] r__65;
  wire [22:0] r__64;
  wire [22:0] r__63;
  wire [22:0] r__62;
  wire [22:0] r__61;
  wire [22:0] r__60;
  wire [22:0] r__59;
  wire [22:0] r__58;
  wire [22:0] r__57;
  wire [22:0] r__56;
  wire [22:0] r__55;
  wire [22:0] r__54;
  wire [22:0] r__53;
  wire [22:0] r__52;
  wire [22:0] r__51;
  wire [22:0] r__50;
  wire [22:0] r__49;
  wire [22:0] r__48;
  wire flag_inf;
  wire [22:0] r__47;
  wire p0_data_enable;
  wire lhs_valid_inv;
  wire rhs_valid_inv;
  wire [22:0] q__23;
  wire [23:0] r__45;
  wire [23:0] r__43;
  wire [23:0] r__41;
  wire [23:0] r__39;
  wire [23:0] r__37;
  wire [23:0] r__35;
  wire [23:0] r__33;
  wire [23:0] r__31;
  wire [23:0] r__29;
  wire [23:0] r__27;
  wire [23:0] r__25;
  wire [23:0] r__23;
  wire [23:0] r__21;
  wire [23:0] r__19;
  wire [23:0] r__17;
  wire [23:0] r__15;
  wire [23:0] r__13;
  wire [23:0] r__11;
  wire [23:0] r__9;
  wire [23:0] r__7;
  wire [23:0] r__5;
  wire [23:0] r__3;
  wire [23:0] b_fractionivisor__1;
  wire [8:0] sub_4129;
  wire b_sign;
  wire [22:0] a_fraction;
  wire lhs_valid_load_en;
  wire rhs_valid_load_en;
  wire [22:0] result_significant;
  wire p30_enable;
  wire p29_enable;
  wire p28_enable;
  wire p27_enable;
  wire p26_enable;
  wire p25_enable;
  wire p24_enable;
  wire q__23_squeezed_portion_0_width_1;
  wire [22:0] concat_5457;
  wire uge_5458;
  wire [22:0] concat_5391;
  wire uge_5392;
  wire [22:0] concat_5325;
  wire uge_5326;
  wire [22:0] concat_5259;
  wire uge_5260;
  wire [22:0] concat_5193;
  wire uge_5194;
  wire [22:0] concat_5127;
  wire uge_5128;
  wire [22:0] concat_5061;
  wire uge_5062;
  wire [22:0] concat_4995;
  wire uge_4996;
  wire [22:0] concat_4929;
  wire uge_4930;
  wire [22:0] concat_4863;
  wire uge_4864;
  wire [22:0] concat_4797;
  wire uge_4798;
  wire [22:0] concat_4731;
  wire uge_4732;
  wire [22:0] concat_4665;
  wire uge_4666;
  wire [22:0] concat_4599;
  wire uge_4600;
  wire [22:0] concat_4533;
  wire uge_4534;
  wire [22:0] concat_4467;
  wire uge_4468;
  wire [22:0] concat_4401;
  wire uge_4402;
  wire [22:0] concat_4335;
  wire uge_4336;
  wire [22:0] concat_4269;
  wire uge_4270;
  wire [22:0] concat_4194;
  wire uge_4195;
  wire [7:0] result_exp;
  wire [22:0] concat_4123;
  wire uge_4124;
  wire [8:0] signed_exp_s9;
  wire [22:0] concat_4053;
  wire [22:0] b_fraction;
  wire [7:0] b_bexp;
  wire result_sign;
  wire bit_slice_3967;
  wire bit_slice_3968;
  wire bit_slice_3969;
  wire bit_slice_3970;
  wire bit_slice_3971;
  wire bit_slice_3972;
  wire bit_slice_3973;
  wire bit_slice_3974;
  wire bit_slice_3975;
  wire bit_slice_3976;
  wire bit_slice_3977;
  wire bit_slice_3978;
  wire bit_slice_3979;
  wire bit_slice_3980;
  wire bit_slice_3981;
  wire bit_slice_3982;
  wire bit_slice_3983;
  wire bit_slice_3984;
  wire bit_slice_3985;
  wire bit_slice_3986;
  wire bit_slice_3987;
  wire [7:0] a_bexp;
  wire bit_slice_3989;
  wire bit_slice_3990;
  wire a_sign;
  wire lhs_load_en;
  wire rhs_load_en;
  wire [31:0] sum;
  assign result_valid_inv = ~result_valid_reg;
  assign result_valid_load_en = result_ready | result_valid_inv;
  assign result_load_en = p23_valid & result_valid_load_en;
  assign p24_stage_done = p23_valid & result_load_en;
  assign p24_not_valid = ~p23_valid;
  assign p23_enable = p24_stage_done | p24_not_valid;
  assign p23_data_enable = p23_enable & p22_valid;
  assign p23_not_valid = ~p22_valid;
  assign p22_enable = p23_data_enable | p23_not_valid;
  assign p22_data_enable = p22_enable & p21_valid;
  assign p22_not_valid = ~p21_valid;
  assign p21_enable = p22_data_enable | p22_not_valid;
  assign p21_data_enable = p21_enable & p20_valid;
  assign p21_not_valid = ~p20_valid;
  assign p20_enable = p21_data_enable | p21_not_valid;
  assign p20_data_enable = p20_enable & p19_valid;
  assign p20_not_valid = ~p19_valid;
  assign p19_enable = p20_data_enable | p20_not_valid;
  assign p19_data_enable = p19_enable & p18_valid;
  assign p19_not_valid = ~p18_valid;
  assign p18_enable = p19_data_enable | p19_not_valid;
  assign p18_data_enable = p18_enable & p17_valid;
  assign p18_not_valid = ~p17_valid;
  assign p17_enable = p18_data_enable | p18_not_valid;
  assign p17_data_enable = p17_enable & p16_valid;
  assign p17_not_valid = ~p16_valid;
  assign p16_enable = p17_data_enable | p17_not_valid;
  assign p16_data_enable = p16_enable & p15_valid;
  assign p16_not_valid = ~p15_valid;
  assign p15_enable = p16_data_enable | p16_not_valid;
  assign p15_data_enable = p15_enable & p14_valid;
  assign p15_not_valid = ~p14_valid;
  assign p14_enable = p15_data_enable | p15_not_valid;
  assign p14_data_enable = p14_enable & p13_valid;
  assign p14_not_valid = ~p13_valid;
  assign p13_enable = p14_data_enable | p14_not_valid;
  assign p13_data_enable = p13_enable & p12_valid;
  assign p13_not_valid = ~p12_valid;
  assign p12_enable = p13_data_enable | p13_not_valid;
  assign p12_data_enable = p12_enable & p11_valid;
  assign p12_not_valid = ~p11_valid;
  assign p11_enable = p12_data_enable | p12_not_valid;
  assign p11_data_enable = p11_enable & p10_valid;
  assign p11_not_valid = ~p10_valid;
  assign p10_enable = p11_data_enable | p11_not_valid;
  assign p10_data_enable = p10_enable & p9_valid;
  assign p10_not_valid = ~p9_valid;
  assign p9_enable = p10_data_enable | p10_not_valid;
  assign p9_data_enable = p9_enable & p8_valid;
  assign p9_not_valid = ~p8_valid;
  assign p8_enable = p9_data_enable | p9_not_valid;
  assign p8_data_enable = p8_enable & p7_valid;
  assign p8_not_valid = ~p7_valid;
  assign p7_enable = p8_data_enable | p8_not_valid;
  assign p7_data_enable = p7_enable & p6_valid;
  assign p7_not_valid = ~p6_valid;
  assign p6_enable = p7_data_enable | p7_not_valid;
  assign p6_data_enable = p6_enable & p5_valid;
  assign p6_not_valid = ~p5_valid;
  assign p5_enable = p6_data_enable | p6_not_valid;
  assign p5_data_enable = p5_enable & p4_valid;
  assign p5_not_valid = ~p4_valid;
  assign p4_enable = p5_data_enable | p5_not_valid;
  assign p4_data_enable = p4_enable & p3_valid;
  assign p4_not_valid = ~p3_valid;
  assign p3_enable = p4_data_enable | p4_not_valid;
  assign p3_data_enable = p3_enable & p2_valid;
  assign p3_not_valid = ~p2_valid;
  assign p2_enable = p3_data_enable | p3_not_valid;
  assign p2_data_enable = p2_enable & p1_valid;
  assign p2_not_valid = ~p1_valid;
  assign p1_enable = p2_data_enable | p2_not_valid;
  assign p1_stage_done = p0_valid & rhs_valid_reg;
  assign p1_data_enable = p1_enable & p1_stage_done;
  assign p1_not_valid = ~p0_valid;
  assign sub_5519 = p22_concat_5457 - p22_b_fraction;
  assign sub_5453 = p21_concat_5391 - p21_b_fraction;
  assign sub_5387 = p20_concat_5325 - p20_b_fraction;
  assign sub_5321 = p19_concat_5259 - p19_b_fraction;
  assign sub_5255 = p18_concat_5193 - p18_b_fraction;
  assign sub_5189 = p17_concat_5127 - p17_b_fraction;
  assign sub_5123 = p16_concat_5061 - p16_b_fraction;
  assign sub_5057 = p15_concat_4995 - p15_b_fraction;
  assign sub_4991 = p14_concat_4929 - p14_b_fraction;
  assign sub_4925 = p13_concat_4863 - p13_b_fraction;
  assign sub_4859 = p12_concat_4797 - p12_b_fraction;
  assign sub_4793 = p11_concat_4731 - p11_b_fraction;
  assign sub_4727 = p10_concat_4665 - p10_b_fraction;
  assign sub_4661 = p9_concat_4599 - p9_b_fraction;
  assign sub_4595 = p8_concat_4533 - p8_b_fraction;
  assign sub_4529 = p7_concat_4467 - p7_b_fraction;
  assign sub_4463 = p6_concat_4401 - p6_b_fraction;
  assign sub_4397 = p5_concat_4335 - p5_b_fraction;
  assign sub_4331 = p4_concat_4269 - p4_b_fraction;
  assign sub_4265 = p3_concat_4194 - p3_b_fraction;
  assign sub_4190 = p2_concat_4123 - p2_b_fraction;
  assign flag_zero = p2_signed_exp_s9[8];
  assign uge_4116 = p1_concat_4053 >= p1_b_fraction;
  assign sub_4117 = p1_concat_4053 - p1_b_fraction;
  assign p0_enable = p1_data_enable | p1_not_valid;
  assign r__68 = p22_uge_5458 ? sub_5519 : p22_concat_5457;
  assign r__67 = p21_uge_5392 ? sub_5453 : p21_concat_5391;
  assign r__66 = p20_uge_5326 ? sub_5387 : p20_concat_5325;
  assign r__65 = p19_uge_5260 ? sub_5321 : p19_concat_5259;
  assign r__64 = p18_uge_5194 ? sub_5255 : p18_concat_5193;
  assign r__63 = p17_uge_5128 ? sub_5189 : p17_concat_5127;
  assign r__62 = p16_uge_5062 ? sub_5123 : p16_concat_5061;
  assign r__61 = p15_uge_4996 ? sub_5057 : p15_concat_4995;
  assign r__60 = p14_uge_4930 ? sub_4991 : p14_concat_4929;
  assign r__59 = p13_uge_4864 ? sub_4925 : p13_concat_4863;
  assign r__58 = p12_uge_4798 ? sub_4859 : p12_concat_4797;
  assign r__57 = p11_uge_4732 ? sub_4793 : p11_concat_4731;
  assign r__56 = p10_uge_4666 ? sub_4727 : p10_concat_4665;
  assign r__55 = p9_uge_4600 ? sub_4661 : p9_concat_4599;
  assign r__54 = p8_uge_4534 ? sub_4595 : p8_concat_4533;
  assign r__53 = p7_uge_4468 ? sub_4529 : p7_concat_4467;
  assign r__52 = p6_uge_4402 ? sub_4463 : p6_concat_4401;
  assign r__51 = p5_uge_4336 ? sub_4397 : p5_concat_4335;
  assign r__50 = p4_uge_4270 ? sub_4331 : p4_concat_4269;
  assign r__49 = p3_uge_4195 ? sub_4265 : p3_concat_4194;
  assign r__48 = p2_uge_4124 ? sub_4190 : p2_concat_4123;
  assign flag_inf = $signed(p2_signed_exp_s9) > $signed(9'h0fe);
  assign r__47 = uge_4116 ? sub_4117 : p1_concat_4053;
  assign p0_data_enable = p0_enable & lhs_valid_reg;
  assign lhs_valid_inv = ~lhs_valid_reg;
  assign rhs_valid_inv = ~rhs_valid_reg;
  assign q__23 = {p23_uge_4116, p23_uge_4124, p23_uge_4195, p23_uge_4270, p23_uge_4336, p23_uge_4402, p23_uge_4468, p23_uge_4534, p23_uge_4600, p23_uge_4666, p23_uge_4732, p23_uge_4798, p23_uge_4864, p23_uge_4930, p23_uge_4996, p23_uge_5062, p23_uge_5128, p23_uge_5194, p23_uge_5260, p23_uge_5326, p23_uge_5392, p23_uge_5458, p23_q__23_squeezed_portion_0_width_1};
  assign r__45 = {r__68, p22_bit_slice_3990};
  assign r__43 = {r__67, p21_bit_slice_3989};
  assign r__41 = {r__66, p20_bit_slice_3987};
  assign r__39 = {r__65, p19_bit_slice_3986};
  assign r__37 = {r__64, p18_bit_slice_3985};
  assign r__35 = {r__63, p17_bit_slice_3984};
  assign r__33 = {r__62, p16_bit_slice_3983};
  assign r__31 = {r__61, p15_bit_slice_3982};
  assign r__29 = {r__60, p14_bit_slice_3981};
  assign r__27 = {r__59, p13_bit_slice_3980};
  assign r__25 = {r__58, p12_bit_slice_3979};
  assign r__23 = {r__57, p11_bit_slice_3978};
  assign r__21 = {r__56, p10_bit_slice_3977};
  assign r__19 = {r__55, p9_bit_slice_3976};
  assign r__17 = {r__54, p8_bit_slice_3975};
  assign r__15 = {r__53, p7_bit_slice_3974};
  assign r__13 = {r__52, p6_bit_slice_3973};
  assign r__11 = {r__51, p5_bit_slice_3972};
  assign r__9 = {r__50, p4_bit_slice_3971};
  assign r__7 = {r__49, p3_bit_slice_3970};
  assign r__5 = {r__48, p2_bit_slice_3969};
  assign r__3 = {r__47, p1_bit_slice_3968};
  assign b_fractionivisor__1 = {1'h0, p1_b_fraction};
  assign sub_4129 = {1'h0, p1_a_bexp} - {1'h0, p1_b_bexp};
  assign b_sign = rhs_reg[31:31];
  assign a_fraction = lhs_reg[22:0];
  assign lhs_valid_load_en = p0_data_enable | lhs_valid_inv;
  assign rhs_valid_load_en = p1_data_enable | rhs_valid_inv;
  assign result_significant = p23_flag_zero ? 23'h00_0001 : q__23;
  assign p30_enable = 1'h1;
  assign p29_enable = 1'h1;
  assign p28_enable = 1'h1;
  assign p27_enable = 1'h1;
  assign p26_enable = 1'h1;
  assign p25_enable = 1'h1;
  assign p24_enable = 1'h1;
  assign q__23_squeezed_portion_0_width_1 = r__45 >= p22_b_fractionivisor__1;
  assign concat_5457 = {r__67[21:0], p21_bit_slice_3989};
  assign uge_5458 = r__43 >= p21_b_fractionivisor__1;
  assign concat_5391 = {r__66[21:0], p20_bit_slice_3987};
  assign uge_5392 = r__41 >= p20_b_fractionivisor__1;
  assign concat_5325 = {r__65[21:0], p19_bit_slice_3986};
  assign uge_5326 = r__39 >= p19_b_fractionivisor__1;
  assign concat_5259 = {r__64[21:0], p18_bit_slice_3985};
  assign uge_5260 = r__37 >= p18_b_fractionivisor__1;
  assign concat_5193 = {r__63[21:0], p17_bit_slice_3984};
  assign uge_5194 = r__35 >= p17_b_fractionivisor__1;
  assign concat_5127 = {r__62[21:0], p16_bit_slice_3983};
  assign uge_5128 = r__33 >= p16_b_fractionivisor__1;
  assign concat_5061 = {r__61[21:0], p15_bit_slice_3982};
  assign uge_5062 = r__31 >= p15_b_fractionivisor__1;
  assign concat_4995 = {r__60[21:0], p14_bit_slice_3981};
  assign uge_4996 = r__29 >= p14_b_fractionivisor__1;
  assign concat_4929 = {r__59[21:0], p13_bit_slice_3980};
  assign uge_4930 = r__27 >= p13_b_fractionivisor__1;
  assign concat_4863 = {r__58[21:0], p12_bit_slice_3979};
  assign uge_4864 = r__25 >= p12_b_fractionivisor__1;
  assign concat_4797 = {r__57[21:0], p11_bit_slice_3978};
  assign uge_4798 = r__23 >= p11_b_fractionivisor__1;
  assign concat_4731 = {r__56[21:0], p10_bit_slice_3977};
  assign uge_4732 = r__21 >= p10_b_fractionivisor__1;
  assign concat_4665 = {r__55[21:0], p9_bit_slice_3976};
  assign uge_4666 = r__19 >= p9_b_fractionivisor__1;
  assign concat_4599 = {r__54[21:0], p8_bit_slice_3975};
  assign uge_4600 = r__17 >= p8_b_fractionivisor__1;
  assign concat_4533 = {r__53[21:0], p7_bit_slice_3974};
  assign uge_4534 = r__15 >= p7_b_fractionivisor__1;
  assign concat_4467 = {r__52[21:0], p6_bit_slice_3973};
  assign uge_4468 = r__13 >= p6_b_fractionivisor__1;
  assign concat_4401 = {r__51[21:0], p5_bit_slice_3972};
  assign uge_4402 = r__11 >= p5_b_fractionivisor__1;
  assign concat_4335 = {r__50[21:0], p4_bit_slice_3971};
  assign uge_4336 = r__9 >= p4_b_fractionivisor__1;
  assign concat_4269 = {r__49[21:0], p3_bit_slice_3970};
  assign uge_4270 = r__7 >= p3_b_fractionivisor__1;
  assign concat_4194 = {r__48[21:0], p2_bit_slice_3969};
  assign uge_4195 = r__5 >= p2_b_fractionivisor__1;
  assign result_exp = (flag_inf ? 8'hff : p2_signed_exp_s9[7:0]) & {8{~flag_zero}};
  assign concat_4123 = {r__47[21:0], p1_bit_slice_3968};
  assign uge_4124 = r__3 >= b_fractionivisor__1;
  assign signed_exp_s9 = sub_4129 + 9'h07f;
  assign concat_4053 = {22'h00_0000, p0_bit_slice_3967};
  assign b_fraction = rhs_reg[22:0];
  assign b_bexp = rhs_reg[30:23];
  assign result_sign = p0_a_sign ^ b_sign;
  assign bit_slice_3967 = a_fraction[22];
  assign bit_slice_3968 = a_fraction[21];
  assign bit_slice_3969 = a_fraction[20];
  assign bit_slice_3970 = a_fraction[19];
  assign bit_slice_3971 = a_fraction[18];
  assign bit_slice_3972 = a_fraction[17];
  assign bit_slice_3973 = a_fraction[16];
  assign bit_slice_3974 = a_fraction[15];
  assign bit_slice_3975 = a_fraction[14];
  assign bit_slice_3976 = a_fraction[13];
  assign bit_slice_3977 = a_fraction[12];
  assign bit_slice_3978 = a_fraction[11];
  assign bit_slice_3979 = a_fraction[10];
  assign bit_slice_3980 = a_fraction[9];
  assign bit_slice_3981 = a_fraction[8];
  assign bit_slice_3982 = a_fraction[7];
  assign bit_slice_3983 = a_fraction[6];
  assign bit_slice_3984 = a_fraction[5];
  assign bit_slice_3985 = a_fraction[4];
  assign bit_slice_3986 = a_fraction[3];
  assign bit_slice_3987 = a_fraction[2];
  assign a_bexp = lhs_reg[30:23];
  assign bit_slice_3989 = a_fraction[1];
  assign bit_slice_3990 = a_fraction[0];
  assign a_sign = lhs_reg[31:31];
  assign lhs_load_en = lhs_valid & lhs_valid_load_en;
  assign rhs_load_en = rhs_valid & rhs_valid_load_en;
  assign sum = {p23_result_sign, p23_result_exp, result_significant};
  always @ (posedge clk) begin
    if (rst) begin
      p0_bit_slice_3967 <= 1'h0;
      p0_bit_slice_3968 <= 1'h0;
      p0_bit_slice_3969 <= 1'h0;
      p0_bit_slice_3970 <= 1'h0;
      p0_bit_slice_3971 <= 1'h0;
      p0_bit_slice_3972 <= 1'h0;
      p0_bit_slice_3973 <= 1'h0;
      p0_bit_slice_3974 <= 1'h0;
      p0_bit_slice_3975 <= 1'h0;
      p0_bit_slice_3976 <= 1'h0;
      p0_bit_slice_3977 <= 1'h0;
      p0_bit_slice_3978 <= 1'h0;
      p0_bit_slice_3979 <= 1'h0;
      p0_bit_slice_3980 <= 1'h0;
      p0_bit_slice_3981 <= 1'h0;
      p0_bit_slice_3982 <= 1'h0;
      p0_bit_slice_3983 <= 1'h0;
      p0_bit_slice_3984 <= 1'h0;
      p0_bit_slice_3985 <= 1'h0;
      p0_bit_slice_3986 <= 1'h0;
      p0_bit_slice_3987 <= 1'h0;
      p0_a_bexp <= 8'h00;
      p0_bit_slice_3989 <= 1'h0;
      p0_bit_slice_3990 <= 1'h0;
      p0_a_sign <= 1'h0;
      p1_concat_4053 <= 23'h00_0000;
      p1_b_fraction <= 23'h00_0000;
      p1_bit_slice_3968 <= 1'h0;
      p1_bit_slice_3969 <= 1'h0;
      p1_bit_slice_3970 <= 1'h0;
      p1_bit_slice_3971 <= 1'h0;
      p1_bit_slice_3972 <= 1'h0;
      p1_bit_slice_3973 <= 1'h0;
      p1_bit_slice_3974 <= 1'h0;
      p1_bit_slice_3975 <= 1'h0;
      p1_bit_slice_3976 <= 1'h0;
      p1_bit_slice_3977 <= 1'h0;
      p1_bit_slice_3978 <= 1'h0;
      p1_bit_slice_3979 <= 1'h0;
      p1_bit_slice_3980 <= 1'h0;
      p1_bit_slice_3981 <= 1'h0;
      p1_bit_slice_3982 <= 1'h0;
      p1_bit_slice_3983 <= 1'h0;
      p1_bit_slice_3984 <= 1'h0;
      p1_bit_slice_3985 <= 1'h0;
      p1_bit_slice_3986 <= 1'h0;
      p1_bit_slice_3987 <= 1'h0;
      p1_a_bexp <= 8'h00;
      p1_b_bexp <= 8'h00;
      p1_bit_slice_3989 <= 1'h0;
      p1_bit_slice_3990 <= 1'h0;
      p1_result_sign <= 1'h0;
      p2_b_fraction <= 23'h00_0000;
      p2_uge_4116 <= 1'h0;
      p2_b_fractionivisor__1 <= 24'h00_0000;
      p2_concat_4123 <= 23'h00_0000;
      p2_uge_4124 <= 1'h0;
      p2_bit_slice_3969 <= 1'h0;
      p2_bit_slice_3970 <= 1'h0;
      p2_bit_slice_3971 <= 1'h0;
      p2_bit_slice_3972 <= 1'h0;
      p2_bit_slice_3973 <= 1'h0;
      p2_bit_slice_3974 <= 1'h0;
      p2_bit_slice_3975 <= 1'h0;
      p2_bit_slice_3976 <= 1'h0;
      p2_bit_slice_3977 <= 1'h0;
      p2_bit_slice_3978 <= 1'h0;
      p2_bit_slice_3979 <= 1'h0;
      p2_bit_slice_3980 <= 1'h0;
      p2_bit_slice_3981 <= 1'h0;
      p2_bit_slice_3982 <= 1'h0;
      p2_bit_slice_3983 <= 1'h0;
      p2_bit_slice_3984 <= 1'h0;
      p2_bit_slice_3985 <= 1'h0;
      p2_bit_slice_3986 <= 1'h0;
      p2_bit_slice_3987 <= 1'h0;
      p2_bit_slice_3989 <= 1'h0;
      p2_signed_exp_s9 <= 9'h000;
      p2_bit_slice_3990 <= 1'h0;
      p2_result_sign <= 1'h0;
      p3_b_fraction <= 23'h00_0000;
      p3_uge_4116 <= 1'h0;
      p3_b_fractionivisor__1 <= 24'h00_0000;
      p3_uge_4124 <= 1'h0;
      p3_concat_4194 <= 23'h00_0000;
      p3_uge_4195 <= 1'h0;
      p3_bit_slice_3970 <= 1'h0;
      p3_bit_slice_3971 <= 1'h0;
      p3_bit_slice_3972 <= 1'h0;
      p3_bit_slice_3973 <= 1'h0;
      p3_bit_slice_3974 <= 1'h0;
      p3_bit_slice_3975 <= 1'h0;
      p3_bit_slice_3976 <= 1'h0;
      p3_bit_slice_3977 <= 1'h0;
      p3_bit_slice_3978 <= 1'h0;
      p3_bit_slice_3979 <= 1'h0;
      p3_bit_slice_3980 <= 1'h0;
      p3_bit_slice_3981 <= 1'h0;
      p3_bit_slice_3982 <= 1'h0;
      p3_bit_slice_3983 <= 1'h0;
      p3_bit_slice_3984 <= 1'h0;
      p3_bit_slice_3985 <= 1'h0;
      p3_bit_slice_3986 <= 1'h0;
      p3_bit_slice_3987 <= 1'h0;
      p3_bit_slice_3989 <= 1'h0;
      p3_bit_slice_3990 <= 1'h0;
      p3_flag_zero <= 1'h0;
      p3_result_sign <= 1'h0;
      p3_result_exp <= 8'h00;
      p4_b_fraction <= 23'h00_0000;
      p4_uge_4116 <= 1'h0;
      p4_b_fractionivisor__1 <= 24'h00_0000;
      p4_uge_4124 <= 1'h0;
      p4_uge_4195 <= 1'h0;
      p4_concat_4269 <= 23'h00_0000;
      p4_uge_4270 <= 1'h0;
      p4_bit_slice_3971 <= 1'h0;
      p4_bit_slice_3972 <= 1'h0;
      p4_bit_slice_3973 <= 1'h0;
      p4_bit_slice_3974 <= 1'h0;
      p4_bit_slice_3975 <= 1'h0;
      p4_bit_slice_3976 <= 1'h0;
      p4_bit_slice_3977 <= 1'h0;
      p4_bit_slice_3978 <= 1'h0;
      p4_bit_slice_3979 <= 1'h0;
      p4_bit_slice_3980 <= 1'h0;
      p4_bit_slice_3981 <= 1'h0;
      p4_bit_slice_3982 <= 1'h0;
      p4_bit_slice_3983 <= 1'h0;
      p4_bit_slice_3984 <= 1'h0;
      p4_bit_slice_3985 <= 1'h0;
      p4_bit_slice_3986 <= 1'h0;
      p4_bit_slice_3987 <= 1'h0;
      p4_bit_slice_3989 <= 1'h0;
      p4_bit_slice_3990 <= 1'h0;
      p4_flag_zero <= 1'h0;
      p4_result_sign <= 1'h0;
      p4_result_exp <= 8'h00;
      p5_b_fraction <= 23'h00_0000;
      p5_uge_4116 <= 1'h0;
      p5_b_fractionivisor__1 <= 24'h00_0000;
      p5_uge_4124 <= 1'h0;
      p5_uge_4195 <= 1'h0;
      p5_uge_4270 <= 1'h0;
      p5_concat_4335 <= 23'h00_0000;
      p5_uge_4336 <= 1'h0;
      p5_bit_slice_3972 <= 1'h0;
      p5_bit_slice_3973 <= 1'h0;
      p5_bit_slice_3974 <= 1'h0;
      p5_bit_slice_3975 <= 1'h0;
      p5_bit_slice_3976 <= 1'h0;
      p5_bit_slice_3977 <= 1'h0;
      p5_bit_slice_3978 <= 1'h0;
      p5_bit_slice_3979 <= 1'h0;
      p5_bit_slice_3980 <= 1'h0;
      p5_bit_slice_3981 <= 1'h0;
      p5_bit_slice_3982 <= 1'h0;
      p5_bit_slice_3983 <= 1'h0;
      p5_bit_slice_3984 <= 1'h0;
      p5_bit_slice_3985 <= 1'h0;
      p5_bit_slice_3986 <= 1'h0;
      p5_bit_slice_3987 <= 1'h0;
      p5_bit_slice_3989 <= 1'h0;
      p5_bit_slice_3990 <= 1'h0;
      p5_flag_zero <= 1'h0;
      p5_result_sign <= 1'h0;
      p5_result_exp <= 8'h00;
      p6_b_fraction <= 23'h00_0000;
      p6_uge_4116 <= 1'h0;
      p6_b_fractionivisor__1 <= 24'h00_0000;
      p6_uge_4124 <= 1'h0;
      p6_uge_4195 <= 1'h0;
      p6_uge_4270 <= 1'h0;
      p6_uge_4336 <= 1'h0;
      p6_concat_4401 <= 23'h00_0000;
      p6_uge_4402 <= 1'h0;
      p6_bit_slice_3973 <= 1'h0;
      p6_bit_slice_3974 <= 1'h0;
      p6_bit_slice_3975 <= 1'h0;
      p6_bit_slice_3976 <= 1'h0;
      p6_bit_slice_3977 <= 1'h0;
      p6_bit_slice_3978 <= 1'h0;
      p6_bit_slice_3979 <= 1'h0;
      p6_bit_slice_3980 <= 1'h0;
      p6_bit_slice_3981 <= 1'h0;
      p6_bit_slice_3982 <= 1'h0;
      p6_bit_slice_3983 <= 1'h0;
      p6_bit_slice_3984 <= 1'h0;
      p6_bit_slice_3985 <= 1'h0;
      p6_bit_slice_3986 <= 1'h0;
      p6_bit_slice_3987 <= 1'h0;
      p6_bit_slice_3989 <= 1'h0;
      p6_bit_slice_3990 <= 1'h0;
      p6_flag_zero <= 1'h0;
      p6_result_sign <= 1'h0;
      p6_result_exp <= 8'h00;
      p7_b_fraction <= 23'h00_0000;
      p7_uge_4116 <= 1'h0;
      p7_b_fractionivisor__1 <= 24'h00_0000;
      p7_uge_4124 <= 1'h0;
      p7_uge_4195 <= 1'h0;
      p7_uge_4270 <= 1'h0;
      p7_uge_4336 <= 1'h0;
      p7_uge_4402 <= 1'h0;
      p7_concat_4467 <= 23'h00_0000;
      p7_uge_4468 <= 1'h0;
      p7_bit_slice_3974 <= 1'h0;
      p7_bit_slice_3975 <= 1'h0;
      p7_bit_slice_3976 <= 1'h0;
      p7_bit_slice_3977 <= 1'h0;
      p7_bit_slice_3978 <= 1'h0;
      p7_bit_slice_3979 <= 1'h0;
      p7_bit_slice_3980 <= 1'h0;
      p7_bit_slice_3981 <= 1'h0;
      p7_bit_slice_3982 <= 1'h0;
      p7_bit_slice_3983 <= 1'h0;
      p7_bit_slice_3984 <= 1'h0;
      p7_bit_slice_3985 <= 1'h0;
      p7_bit_slice_3986 <= 1'h0;
      p7_bit_slice_3987 <= 1'h0;
      p7_bit_slice_3989 <= 1'h0;
      p7_bit_slice_3990 <= 1'h0;
      p7_flag_zero <= 1'h0;
      p7_result_sign <= 1'h0;
      p7_result_exp <= 8'h00;
      p8_b_fraction <= 23'h00_0000;
      p8_uge_4116 <= 1'h0;
      p8_b_fractionivisor__1 <= 24'h00_0000;
      p8_uge_4124 <= 1'h0;
      p8_uge_4195 <= 1'h0;
      p8_uge_4270 <= 1'h0;
      p8_uge_4336 <= 1'h0;
      p8_uge_4402 <= 1'h0;
      p8_uge_4468 <= 1'h0;
      p8_concat_4533 <= 23'h00_0000;
      p8_uge_4534 <= 1'h0;
      p8_bit_slice_3975 <= 1'h0;
      p8_bit_slice_3976 <= 1'h0;
      p8_bit_slice_3977 <= 1'h0;
      p8_bit_slice_3978 <= 1'h0;
      p8_bit_slice_3979 <= 1'h0;
      p8_bit_slice_3980 <= 1'h0;
      p8_bit_slice_3981 <= 1'h0;
      p8_bit_slice_3982 <= 1'h0;
      p8_bit_slice_3983 <= 1'h0;
      p8_bit_slice_3984 <= 1'h0;
      p8_bit_slice_3985 <= 1'h0;
      p8_bit_slice_3986 <= 1'h0;
      p8_bit_slice_3987 <= 1'h0;
      p8_bit_slice_3989 <= 1'h0;
      p8_bit_slice_3990 <= 1'h0;
      p8_flag_zero <= 1'h0;
      p8_result_sign <= 1'h0;
      p8_result_exp <= 8'h00;
      p9_b_fraction <= 23'h00_0000;
      p9_uge_4116 <= 1'h0;
      p9_b_fractionivisor__1 <= 24'h00_0000;
      p9_uge_4124 <= 1'h0;
      p9_uge_4195 <= 1'h0;
      p9_uge_4270 <= 1'h0;
      p9_uge_4336 <= 1'h0;
      p9_uge_4402 <= 1'h0;
      p9_uge_4468 <= 1'h0;
      p9_uge_4534 <= 1'h0;
      p9_concat_4599 <= 23'h00_0000;
      p9_uge_4600 <= 1'h0;
      p9_bit_slice_3976 <= 1'h0;
      p9_bit_slice_3977 <= 1'h0;
      p9_bit_slice_3978 <= 1'h0;
      p9_bit_slice_3979 <= 1'h0;
      p9_bit_slice_3980 <= 1'h0;
      p9_bit_slice_3981 <= 1'h0;
      p9_bit_slice_3982 <= 1'h0;
      p9_bit_slice_3983 <= 1'h0;
      p9_bit_slice_3984 <= 1'h0;
      p9_bit_slice_3985 <= 1'h0;
      p9_bit_slice_3986 <= 1'h0;
      p9_bit_slice_3987 <= 1'h0;
      p9_bit_slice_3989 <= 1'h0;
      p9_bit_slice_3990 <= 1'h0;
      p9_flag_zero <= 1'h0;
      p9_result_sign <= 1'h0;
      p9_result_exp <= 8'h00;
      p10_b_fraction <= 23'h00_0000;
      p10_uge_4116 <= 1'h0;
      p10_b_fractionivisor__1 <= 24'h00_0000;
      p10_uge_4124 <= 1'h0;
      p10_uge_4195 <= 1'h0;
      p10_uge_4270 <= 1'h0;
      p10_uge_4336 <= 1'h0;
      p10_uge_4402 <= 1'h0;
      p10_uge_4468 <= 1'h0;
      p10_uge_4534 <= 1'h0;
      p10_uge_4600 <= 1'h0;
      p10_concat_4665 <= 23'h00_0000;
      p10_uge_4666 <= 1'h0;
      p10_bit_slice_3977 <= 1'h0;
      p10_bit_slice_3978 <= 1'h0;
      p10_bit_slice_3979 <= 1'h0;
      p10_bit_slice_3980 <= 1'h0;
      p10_bit_slice_3981 <= 1'h0;
      p10_bit_slice_3982 <= 1'h0;
      p10_bit_slice_3983 <= 1'h0;
      p10_bit_slice_3984 <= 1'h0;
      p10_bit_slice_3985 <= 1'h0;
      p10_bit_slice_3986 <= 1'h0;
      p10_bit_slice_3987 <= 1'h0;
      p10_bit_slice_3989 <= 1'h0;
      p10_bit_slice_3990 <= 1'h0;
      p10_flag_zero <= 1'h0;
      p10_result_sign <= 1'h0;
      p10_result_exp <= 8'h00;
      p11_b_fraction <= 23'h00_0000;
      p11_uge_4116 <= 1'h0;
      p11_b_fractionivisor__1 <= 24'h00_0000;
      p11_uge_4124 <= 1'h0;
      p11_uge_4195 <= 1'h0;
      p11_uge_4270 <= 1'h0;
      p11_uge_4336 <= 1'h0;
      p11_uge_4402 <= 1'h0;
      p11_uge_4468 <= 1'h0;
      p11_uge_4534 <= 1'h0;
      p11_uge_4600 <= 1'h0;
      p11_uge_4666 <= 1'h0;
      p11_concat_4731 <= 23'h00_0000;
      p11_uge_4732 <= 1'h0;
      p11_bit_slice_3978 <= 1'h0;
      p11_bit_slice_3979 <= 1'h0;
      p11_bit_slice_3980 <= 1'h0;
      p11_bit_slice_3981 <= 1'h0;
      p11_bit_slice_3982 <= 1'h0;
      p11_bit_slice_3983 <= 1'h0;
      p11_bit_slice_3984 <= 1'h0;
      p11_bit_slice_3985 <= 1'h0;
      p11_bit_slice_3986 <= 1'h0;
      p11_bit_slice_3987 <= 1'h0;
      p11_bit_slice_3989 <= 1'h0;
      p11_bit_slice_3990 <= 1'h0;
      p11_flag_zero <= 1'h0;
      p11_result_sign <= 1'h0;
      p11_result_exp <= 8'h00;
      p12_b_fraction <= 23'h00_0000;
      p12_uge_4116 <= 1'h0;
      p12_b_fractionivisor__1 <= 24'h00_0000;
      p12_uge_4124 <= 1'h0;
      p12_uge_4195 <= 1'h0;
      p12_uge_4270 <= 1'h0;
      p12_uge_4336 <= 1'h0;
      p12_uge_4402 <= 1'h0;
      p12_uge_4468 <= 1'h0;
      p12_uge_4534 <= 1'h0;
      p12_uge_4600 <= 1'h0;
      p12_uge_4666 <= 1'h0;
      p12_uge_4732 <= 1'h0;
      p12_concat_4797 <= 23'h00_0000;
      p12_uge_4798 <= 1'h0;
      p12_bit_slice_3979 <= 1'h0;
      p12_bit_slice_3980 <= 1'h0;
      p12_bit_slice_3981 <= 1'h0;
      p12_bit_slice_3982 <= 1'h0;
      p12_bit_slice_3983 <= 1'h0;
      p12_bit_slice_3984 <= 1'h0;
      p12_bit_slice_3985 <= 1'h0;
      p12_bit_slice_3986 <= 1'h0;
      p12_bit_slice_3987 <= 1'h0;
      p12_bit_slice_3989 <= 1'h0;
      p12_bit_slice_3990 <= 1'h0;
      p12_flag_zero <= 1'h0;
      p12_result_sign <= 1'h0;
      p12_result_exp <= 8'h00;
      p13_b_fraction <= 23'h00_0000;
      p13_uge_4116 <= 1'h0;
      p13_b_fractionivisor__1 <= 24'h00_0000;
      p13_uge_4124 <= 1'h0;
      p13_uge_4195 <= 1'h0;
      p13_uge_4270 <= 1'h0;
      p13_uge_4336 <= 1'h0;
      p13_uge_4402 <= 1'h0;
      p13_uge_4468 <= 1'h0;
      p13_uge_4534 <= 1'h0;
      p13_uge_4600 <= 1'h0;
      p13_uge_4666 <= 1'h0;
      p13_uge_4732 <= 1'h0;
      p13_uge_4798 <= 1'h0;
      p13_concat_4863 <= 23'h00_0000;
      p13_uge_4864 <= 1'h0;
      p13_bit_slice_3980 <= 1'h0;
      p13_bit_slice_3981 <= 1'h0;
      p13_bit_slice_3982 <= 1'h0;
      p13_bit_slice_3983 <= 1'h0;
      p13_bit_slice_3984 <= 1'h0;
      p13_bit_slice_3985 <= 1'h0;
      p13_bit_slice_3986 <= 1'h0;
      p13_bit_slice_3987 <= 1'h0;
      p13_bit_slice_3989 <= 1'h0;
      p13_bit_slice_3990 <= 1'h0;
      p13_flag_zero <= 1'h0;
      p13_result_sign <= 1'h0;
      p13_result_exp <= 8'h00;
      p14_b_fraction <= 23'h00_0000;
      p14_uge_4116 <= 1'h0;
      p14_b_fractionivisor__1 <= 24'h00_0000;
      p14_uge_4124 <= 1'h0;
      p14_uge_4195 <= 1'h0;
      p14_uge_4270 <= 1'h0;
      p14_uge_4336 <= 1'h0;
      p14_uge_4402 <= 1'h0;
      p14_uge_4468 <= 1'h0;
      p14_uge_4534 <= 1'h0;
      p14_uge_4600 <= 1'h0;
      p14_uge_4666 <= 1'h0;
      p14_uge_4732 <= 1'h0;
      p14_uge_4798 <= 1'h0;
      p14_uge_4864 <= 1'h0;
      p14_concat_4929 <= 23'h00_0000;
      p14_uge_4930 <= 1'h0;
      p14_bit_slice_3981 <= 1'h0;
      p14_bit_slice_3982 <= 1'h0;
      p14_bit_slice_3983 <= 1'h0;
      p14_bit_slice_3984 <= 1'h0;
      p14_bit_slice_3985 <= 1'h0;
      p14_bit_slice_3986 <= 1'h0;
      p14_bit_slice_3987 <= 1'h0;
      p14_bit_slice_3989 <= 1'h0;
      p14_bit_slice_3990 <= 1'h0;
      p14_flag_zero <= 1'h0;
      p14_result_sign <= 1'h0;
      p14_result_exp <= 8'h00;
      p15_b_fraction <= 23'h00_0000;
      p15_uge_4116 <= 1'h0;
      p15_b_fractionivisor__1 <= 24'h00_0000;
      p15_uge_4124 <= 1'h0;
      p15_uge_4195 <= 1'h0;
      p15_uge_4270 <= 1'h0;
      p15_uge_4336 <= 1'h0;
      p15_uge_4402 <= 1'h0;
      p15_uge_4468 <= 1'h0;
      p15_uge_4534 <= 1'h0;
      p15_uge_4600 <= 1'h0;
      p15_uge_4666 <= 1'h0;
      p15_uge_4732 <= 1'h0;
      p15_uge_4798 <= 1'h0;
      p15_uge_4864 <= 1'h0;
      p15_uge_4930 <= 1'h0;
      p15_concat_4995 <= 23'h00_0000;
      p15_uge_4996 <= 1'h0;
      p15_bit_slice_3982 <= 1'h0;
      p15_bit_slice_3983 <= 1'h0;
      p15_bit_slice_3984 <= 1'h0;
      p15_bit_slice_3985 <= 1'h0;
      p15_bit_slice_3986 <= 1'h0;
      p15_bit_slice_3987 <= 1'h0;
      p15_bit_slice_3989 <= 1'h0;
      p15_bit_slice_3990 <= 1'h0;
      p15_flag_zero <= 1'h0;
      p15_result_sign <= 1'h0;
      p15_result_exp <= 8'h00;
      p16_b_fraction <= 23'h00_0000;
      p16_uge_4116 <= 1'h0;
      p16_b_fractionivisor__1 <= 24'h00_0000;
      p16_uge_4124 <= 1'h0;
      p16_uge_4195 <= 1'h0;
      p16_uge_4270 <= 1'h0;
      p16_uge_4336 <= 1'h0;
      p16_uge_4402 <= 1'h0;
      p16_uge_4468 <= 1'h0;
      p16_uge_4534 <= 1'h0;
      p16_uge_4600 <= 1'h0;
      p16_uge_4666 <= 1'h0;
      p16_uge_4732 <= 1'h0;
      p16_uge_4798 <= 1'h0;
      p16_uge_4864 <= 1'h0;
      p16_uge_4930 <= 1'h0;
      p16_uge_4996 <= 1'h0;
      p16_concat_5061 <= 23'h00_0000;
      p16_uge_5062 <= 1'h0;
      p16_bit_slice_3983 <= 1'h0;
      p16_bit_slice_3984 <= 1'h0;
      p16_bit_slice_3985 <= 1'h0;
      p16_bit_slice_3986 <= 1'h0;
      p16_bit_slice_3987 <= 1'h0;
      p16_bit_slice_3989 <= 1'h0;
      p16_bit_slice_3990 <= 1'h0;
      p16_flag_zero <= 1'h0;
      p16_result_sign <= 1'h0;
      p16_result_exp <= 8'h00;
      p17_b_fraction <= 23'h00_0000;
      p17_uge_4116 <= 1'h0;
      p17_b_fractionivisor__1 <= 24'h00_0000;
      p17_uge_4124 <= 1'h0;
      p17_uge_4195 <= 1'h0;
      p17_uge_4270 <= 1'h0;
      p17_uge_4336 <= 1'h0;
      p17_uge_4402 <= 1'h0;
      p17_uge_4468 <= 1'h0;
      p17_uge_4534 <= 1'h0;
      p17_uge_4600 <= 1'h0;
      p17_uge_4666 <= 1'h0;
      p17_uge_4732 <= 1'h0;
      p17_uge_4798 <= 1'h0;
      p17_uge_4864 <= 1'h0;
      p17_uge_4930 <= 1'h0;
      p17_uge_4996 <= 1'h0;
      p17_uge_5062 <= 1'h0;
      p17_concat_5127 <= 23'h00_0000;
      p17_uge_5128 <= 1'h0;
      p17_bit_slice_3984 <= 1'h0;
      p17_bit_slice_3985 <= 1'h0;
      p17_bit_slice_3986 <= 1'h0;
      p17_bit_slice_3987 <= 1'h0;
      p17_bit_slice_3989 <= 1'h0;
      p17_bit_slice_3990 <= 1'h0;
      p17_flag_zero <= 1'h0;
      p17_result_sign <= 1'h0;
      p17_result_exp <= 8'h00;
      p18_b_fraction <= 23'h00_0000;
      p18_uge_4116 <= 1'h0;
      p18_b_fractionivisor__1 <= 24'h00_0000;
      p18_uge_4124 <= 1'h0;
      p18_uge_4195 <= 1'h0;
      p18_uge_4270 <= 1'h0;
      p18_uge_4336 <= 1'h0;
      p18_uge_4402 <= 1'h0;
      p18_uge_4468 <= 1'h0;
      p18_uge_4534 <= 1'h0;
      p18_uge_4600 <= 1'h0;
      p18_uge_4666 <= 1'h0;
      p18_uge_4732 <= 1'h0;
      p18_uge_4798 <= 1'h0;
      p18_uge_4864 <= 1'h0;
      p18_uge_4930 <= 1'h0;
      p18_uge_4996 <= 1'h0;
      p18_uge_5062 <= 1'h0;
      p18_uge_5128 <= 1'h0;
      p18_concat_5193 <= 23'h00_0000;
      p18_uge_5194 <= 1'h0;
      p18_bit_slice_3985 <= 1'h0;
      p18_bit_slice_3986 <= 1'h0;
      p18_bit_slice_3987 <= 1'h0;
      p18_bit_slice_3989 <= 1'h0;
      p18_bit_slice_3990 <= 1'h0;
      p18_flag_zero <= 1'h0;
      p18_result_sign <= 1'h0;
      p18_result_exp <= 8'h00;
      p19_b_fraction <= 23'h00_0000;
      p19_uge_4116 <= 1'h0;
      p19_b_fractionivisor__1 <= 24'h00_0000;
      p19_uge_4124 <= 1'h0;
      p19_uge_4195 <= 1'h0;
      p19_uge_4270 <= 1'h0;
      p19_uge_4336 <= 1'h0;
      p19_uge_4402 <= 1'h0;
      p19_uge_4468 <= 1'h0;
      p19_uge_4534 <= 1'h0;
      p19_uge_4600 <= 1'h0;
      p19_uge_4666 <= 1'h0;
      p19_uge_4732 <= 1'h0;
      p19_uge_4798 <= 1'h0;
      p19_uge_4864 <= 1'h0;
      p19_uge_4930 <= 1'h0;
      p19_uge_4996 <= 1'h0;
      p19_uge_5062 <= 1'h0;
      p19_uge_5128 <= 1'h0;
      p19_uge_5194 <= 1'h0;
      p19_concat_5259 <= 23'h00_0000;
      p19_uge_5260 <= 1'h0;
      p19_bit_slice_3986 <= 1'h0;
      p19_bit_slice_3987 <= 1'h0;
      p19_bit_slice_3989 <= 1'h0;
      p19_bit_slice_3990 <= 1'h0;
      p19_flag_zero <= 1'h0;
      p19_result_sign <= 1'h0;
      p19_result_exp <= 8'h00;
      p20_b_fraction <= 23'h00_0000;
      p20_uge_4116 <= 1'h0;
      p20_b_fractionivisor__1 <= 24'h00_0000;
      p20_uge_4124 <= 1'h0;
      p20_uge_4195 <= 1'h0;
      p20_uge_4270 <= 1'h0;
      p20_uge_4336 <= 1'h0;
      p20_uge_4402 <= 1'h0;
      p20_uge_4468 <= 1'h0;
      p20_uge_4534 <= 1'h0;
      p20_uge_4600 <= 1'h0;
      p20_uge_4666 <= 1'h0;
      p20_uge_4732 <= 1'h0;
      p20_uge_4798 <= 1'h0;
      p20_uge_4864 <= 1'h0;
      p20_uge_4930 <= 1'h0;
      p20_uge_4996 <= 1'h0;
      p20_uge_5062 <= 1'h0;
      p20_uge_5128 <= 1'h0;
      p20_uge_5194 <= 1'h0;
      p20_uge_5260 <= 1'h0;
      p20_concat_5325 <= 23'h00_0000;
      p20_uge_5326 <= 1'h0;
      p20_bit_slice_3987 <= 1'h0;
      p20_bit_slice_3989 <= 1'h0;
      p20_bit_slice_3990 <= 1'h0;
      p20_flag_zero <= 1'h0;
      p20_result_sign <= 1'h0;
      p20_result_exp <= 8'h00;
      p21_b_fraction <= 23'h00_0000;
      p21_uge_4116 <= 1'h0;
      p21_b_fractionivisor__1 <= 24'h00_0000;
      p21_uge_4124 <= 1'h0;
      p21_uge_4195 <= 1'h0;
      p21_uge_4270 <= 1'h0;
      p21_uge_4336 <= 1'h0;
      p21_uge_4402 <= 1'h0;
      p21_uge_4468 <= 1'h0;
      p21_uge_4534 <= 1'h0;
      p21_uge_4600 <= 1'h0;
      p21_uge_4666 <= 1'h0;
      p21_uge_4732 <= 1'h0;
      p21_uge_4798 <= 1'h0;
      p21_uge_4864 <= 1'h0;
      p21_uge_4930 <= 1'h0;
      p21_uge_4996 <= 1'h0;
      p21_uge_5062 <= 1'h0;
      p21_uge_5128 <= 1'h0;
      p21_uge_5194 <= 1'h0;
      p21_uge_5260 <= 1'h0;
      p21_uge_5326 <= 1'h0;
      p21_concat_5391 <= 23'h00_0000;
      p21_uge_5392 <= 1'h0;
      p21_bit_slice_3989 <= 1'h0;
      p21_bit_slice_3990 <= 1'h0;
      p21_flag_zero <= 1'h0;
      p21_result_sign <= 1'h0;
      p21_result_exp <= 8'h00;
      p22_b_fraction <= 23'h00_0000;
      p22_uge_4116 <= 1'h0;
      p22_b_fractionivisor__1 <= 24'h00_0000;
      p22_uge_4124 <= 1'h0;
      p22_uge_4195 <= 1'h0;
      p22_uge_4270 <= 1'h0;
      p22_uge_4336 <= 1'h0;
      p22_uge_4402 <= 1'h0;
      p22_uge_4468 <= 1'h0;
      p22_uge_4534 <= 1'h0;
      p22_uge_4600 <= 1'h0;
      p22_uge_4666 <= 1'h0;
      p22_uge_4732 <= 1'h0;
      p22_uge_4798 <= 1'h0;
      p22_uge_4864 <= 1'h0;
      p22_uge_4930 <= 1'h0;
      p22_uge_4996 <= 1'h0;
      p22_uge_5062 <= 1'h0;
      p22_uge_5128 <= 1'h0;
      p22_uge_5194 <= 1'h0;
      p22_uge_5260 <= 1'h0;
      p22_uge_5326 <= 1'h0;
      p22_uge_5392 <= 1'h0;
      p22_concat_5457 <= 23'h00_0000;
      p22_uge_5458 <= 1'h0;
      p22_bit_slice_3990 <= 1'h0;
      p22_flag_zero <= 1'h0;
      p22_result_sign <= 1'h0;
      p22_result_exp <= 8'h00;
      p23_uge_4116 <= 1'h0;
      p23_uge_4124 <= 1'h0;
      p23_uge_4195 <= 1'h0;
      p23_uge_4270 <= 1'h0;
      p23_uge_4336 <= 1'h0;
      p23_uge_4402 <= 1'h0;
      p23_uge_4468 <= 1'h0;
      p23_uge_4534 <= 1'h0;
      p23_uge_4600 <= 1'h0;
      p23_uge_4666 <= 1'h0;
      p23_uge_4732 <= 1'h0;
      p23_uge_4798 <= 1'h0;
      p23_uge_4864 <= 1'h0;
      p23_uge_4930 <= 1'h0;
      p23_uge_4996 <= 1'h0;
      p23_uge_5062 <= 1'h0;
      p23_uge_5128 <= 1'h0;
      p23_uge_5194 <= 1'h0;
      p23_uge_5260 <= 1'h0;
      p23_uge_5326 <= 1'h0;
      p23_uge_5392 <= 1'h0;
      p23_uge_5458 <= 1'h0;
      p23_flag_zero <= 1'h0;
      p23_q__23_squeezed_portion_0_width_1 <= 1'h0;
      p23_result_sign <= 1'h0;
      p23_result_exp <= 8'h00;
      p0_valid <= 1'h0;
      p1_valid <= 1'h0;
      p2_valid <= 1'h0;
      p3_valid <= 1'h0;
      p4_valid <= 1'h0;
      p5_valid <= 1'h0;
      p6_valid <= 1'h0;
      p7_valid <= 1'h0;
      p8_valid <= 1'h0;
      p9_valid <= 1'h0;
      p10_valid <= 1'h0;
      p11_valid <= 1'h0;
      p12_valid <= 1'h0;
      p13_valid <= 1'h0;
      p14_valid <= 1'h0;
      p15_valid <= 1'h0;
      p16_valid <= 1'h0;
      p17_valid <= 1'h0;
      p18_valid <= 1'h0;
      p19_valid <= 1'h0;
      p20_valid <= 1'h0;
      p21_valid <= 1'h0;
      p22_valid <= 1'h0;
      p23_valid <= 1'h0;
      p24_valid <= 1'h0;
      p25_valid <= 1'h0;
      p26_valid <= 1'h0;
      p27_valid <= 1'h0;
      p28_valid <= 1'h0;
      p29_valid <= 1'h0;
      p30_valid <= 1'h0;
      lhs_reg <= lhs_reg_init;
      lhs_valid_reg <= 1'h0;
      rhs_reg <= rhs_reg_init;
      rhs_valid_reg <= 1'h0;
      result_reg <= result_reg_init;
      result_valid_reg <= 1'h0;
    end else begin
      p0_bit_slice_3967 <= p0_data_enable ? bit_slice_3967 : p0_bit_slice_3967;
      p0_bit_slice_3968 <= p0_data_enable ? bit_slice_3968 : p0_bit_slice_3968;
      p0_bit_slice_3969 <= p0_data_enable ? bit_slice_3969 : p0_bit_slice_3969;
      p0_bit_slice_3970 <= p0_data_enable ? bit_slice_3970 : p0_bit_slice_3970;
      p0_bit_slice_3971 <= p0_data_enable ? bit_slice_3971 : p0_bit_slice_3971;
      p0_bit_slice_3972 <= p0_data_enable ? bit_slice_3972 : p0_bit_slice_3972;
      p0_bit_slice_3973 <= p0_data_enable ? bit_slice_3973 : p0_bit_slice_3973;
      p0_bit_slice_3974 <= p0_data_enable ? bit_slice_3974 : p0_bit_slice_3974;
      p0_bit_slice_3975 <= p0_data_enable ? bit_slice_3975 : p0_bit_slice_3975;
      p0_bit_slice_3976 <= p0_data_enable ? bit_slice_3976 : p0_bit_slice_3976;
      p0_bit_slice_3977 <= p0_data_enable ? bit_slice_3977 : p0_bit_slice_3977;
      p0_bit_slice_3978 <= p0_data_enable ? bit_slice_3978 : p0_bit_slice_3978;
      p0_bit_slice_3979 <= p0_data_enable ? bit_slice_3979 : p0_bit_slice_3979;
      p0_bit_slice_3980 <= p0_data_enable ? bit_slice_3980 : p0_bit_slice_3980;
      p0_bit_slice_3981 <= p0_data_enable ? bit_slice_3981 : p0_bit_slice_3981;
      p0_bit_slice_3982 <= p0_data_enable ? bit_slice_3982 : p0_bit_slice_3982;
      p0_bit_slice_3983 <= p0_data_enable ? bit_slice_3983 : p0_bit_slice_3983;
      p0_bit_slice_3984 <= p0_data_enable ? bit_slice_3984 : p0_bit_slice_3984;
      p0_bit_slice_3985 <= p0_data_enable ? bit_slice_3985 : p0_bit_slice_3985;
      p0_bit_slice_3986 <= p0_data_enable ? bit_slice_3986 : p0_bit_slice_3986;
      p0_bit_slice_3987 <= p0_data_enable ? bit_slice_3987 : p0_bit_slice_3987;
      p0_a_bexp <= p0_data_enable ? a_bexp : p0_a_bexp;
      p0_bit_slice_3989 <= p0_data_enable ? bit_slice_3989 : p0_bit_slice_3989;
      p0_bit_slice_3990 <= p0_data_enable ? bit_slice_3990 : p0_bit_slice_3990;
      p0_a_sign <= p0_data_enable ? a_sign : p0_a_sign;
      p1_concat_4053 <= p1_data_enable ? concat_4053 : p1_concat_4053;
      p1_b_fraction <= p1_data_enable ? b_fraction : p1_b_fraction;
      p1_bit_slice_3968 <= p1_data_enable ? p0_bit_slice_3968 : p1_bit_slice_3968;
      p1_bit_slice_3969 <= p1_data_enable ? p0_bit_slice_3969 : p1_bit_slice_3969;
      p1_bit_slice_3970 <= p1_data_enable ? p0_bit_slice_3970 : p1_bit_slice_3970;
      p1_bit_slice_3971 <= p1_data_enable ? p0_bit_slice_3971 : p1_bit_slice_3971;
      p1_bit_slice_3972 <= p1_data_enable ? p0_bit_slice_3972 : p1_bit_slice_3972;
      p1_bit_slice_3973 <= p1_data_enable ? p0_bit_slice_3973 : p1_bit_slice_3973;
      p1_bit_slice_3974 <= p1_data_enable ? p0_bit_slice_3974 : p1_bit_slice_3974;
      p1_bit_slice_3975 <= p1_data_enable ? p0_bit_slice_3975 : p1_bit_slice_3975;
      p1_bit_slice_3976 <= p1_data_enable ? p0_bit_slice_3976 : p1_bit_slice_3976;
      p1_bit_slice_3977 <= p1_data_enable ? p0_bit_slice_3977 : p1_bit_slice_3977;
      p1_bit_slice_3978 <= p1_data_enable ? p0_bit_slice_3978 : p1_bit_slice_3978;
      p1_bit_slice_3979 <= p1_data_enable ? p0_bit_slice_3979 : p1_bit_slice_3979;
      p1_bit_slice_3980 <= p1_data_enable ? p0_bit_slice_3980 : p1_bit_slice_3980;
      p1_bit_slice_3981 <= p1_data_enable ? p0_bit_slice_3981 : p1_bit_slice_3981;
      p1_bit_slice_3982 <= p1_data_enable ? p0_bit_slice_3982 : p1_bit_slice_3982;
      p1_bit_slice_3983 <= p1_data_enable ? p0_bit_slice_3983 : p1_bit_slice_3983;
      p1_bit_slice_3984 <= p1_data_enable ? p0_bit_slice_3984 : p1_bit_slice_3984;
      p1_bit_slice_3985 <= p1_data_enable ? p0_bit_slice_3985 : p1_bit_slice_3985;
      p1_bit_slice_3986 <= p1_data_enable ? p0_bit_slice_3986 : p1_bit_slice_3986;
      p1_bit_slice_3987 <= p1_data_enable ? p0_bit_slice_3987 : p1_bit_slice_3987;
      p1_a_bexp <= p1_data_enable ? p0_a_bexp : p1_a_bexp;
      p1_b_bexp <= p1_data_enable ? b_bexp : p1_b_bexp;
      p1_bit_slice_3989 <= p1_data_enable ? p0_bit_slice_3989 : p1_bit_slice_3989;
      p1_bit_slice_3990 <= p1_data_enable ? p0_bit_slice_3990 : p1_bit_slice_3990;
      p1_result_sign <= p1_data_enable ? result_sign : p1_result_sign;
      p2_b_fraction <= p2_data_enable ? p1_b_fraction : p2_b_fraction;
      p2_uge_4116 <= p2_data_enable ? uge_4116 : p2_uge_4116;
      p2_b_fractionivisor__1 <= p2_data_enable ? b_fractionivisor__1 : p2_b_fractionivisor__1;
      p2_concat_4123 <= p2_data_enable ? concat_4123 : p2_concat_4123;
      p2_uge_4124 <= p2_data_enable ? uge_4124 : p2_uge_4124;
      p2_bit_slice_3969 <= p2_data_enable ? p1_bit_slice_3969 : p2_bit_slice_3969;
      p2_bit_slice_3970 <= p2_data_enable ? p1_bit_slice_3970 : p2_bit_slice_3970;
      p2_bit_slice_3971 <= p2_data_enable ? p1_bit_slice_3971 : p2_bit_slice_3971;
      p2_bit_slice_3972 <= p2_data_enable ? p1_bit_slice_3972 : p2_bit_slice_3972;
      p2_bit_slice_3973 <= p2_data_enable ? p1_bit_slice_3973 : p2_bit_slice_3973;
      p2_bit_slice_3974 <= p2_data_enable ? p1_bit_slice_3974 : p2_bit_slice_3974;
      p2_bit_slice_3975 <= p2_data_enable ? p1_bit_slice_3975 : p2_bit_slice_3975;
      p2_bit_slice_3976 <= p2_data_enable ? p1_bit_slice_3976 : p2_bit_slice_3976;
      p2_bit_slice_3977 <= p2_data_enable ? p1_bit_slice_3977 : p2_bit_slice_3977;
      p2_bit_slice_3978 <= p2_data_enable ? p1_bit_slice_3978 : p2_bit_slice_3978;
      p2_bit_slice_3979 <= p2_data_enable ? p1_bit_slice_3979 : p2_bit_slice_3979;
      p2_bit_slice_3980 <= p2_data_enable ? p1_bit_slice_3980 : p2_bit_slice_3980;
      p2_bit_slice_3981 <= p2_data_enable ? p1_bit_slice_3981 : p2_bit_slice_3981;
      p2_bit_slice_3982 <= p2_data_enable ? p1_bit_slice_3982 : p2_bit_slice_3982;
      p2_bit_slice_3983 <= p2_data_enable ? p1_bit_slice_3983 : p2_bit_slice_3983;
      p2_bit_slice_3984 <= p2_data_enable ? p1_bit_slice_3984 : p2_bit_slice_3984;
      p2_bit_slice_3985 <= p2_data_enable ? p1_bit_slice_3985 : p2_bit_slice_3985;
      p2_bit_slice_3986 <= p2_data_enable ? p1_bit_slice_3986 : p2_bit_slice_3986;
      p2_bit_slice_3987 <= p2_data_enable ? p1_bit_slice_3987 : p2_bit_slice_3987;
      p2_bit_slice_3989 <= p2_data_enable ? p1_bit_slice_3989 : p2_bit_slice_3989;
      p2_signed_exp_s9 <= p2_data_enable ? signed_exp_s9 : p2_signed_exp_s9;
      p2_bit_slice_3990 <= p2_data_enable ? p1_bit_slice_3990 : p2_bit_slice_3990;
      p2_result_sign <= p2_data_enable ? p1_result_sign : p2_result_sign;
      p3_b_fraction <= p3_data_enable ? p2_b_fraction : p3_b_fraction;
      p3_uge_4116 <= p3_data_enable ? p2_uge_4116 : p3_uge_4116;
      p3_b_fractionivisor__1 <= p3_data_enable ? p2_b_fractionivisor__1 : p3_b_fractionivisor__1;
      p3_uge_4124 <= p3_data_enable ? p2_uge_4124 : p3_uge_4124;
      p3_concat_4194 <= p3_data_enable ? concat_4194 : p3_concat_4194;
      p3_uge_4195 <= p3_data_enable ? uge_4195 : p3_uge_4195;
      p3_bit_slice_3970 <= p3_data_enable ? p2_bit_slice_3970 : p3_bit_slice_3970;
      p3_bit_slice_3971 <= p3_data_enable ? p2_bit_slice_3971 : p3_bit_slice_3971;
      p3_bit_slice_3972 <= p3_data_enable ? p2_bit_slice_3972 : p3_bit_slice_3972;
      p3_bit_slice_3973 <= p3_data_enable ? p2_bit_slice_3973 : p3_bit_slice_3973;
      p3_bit_slice_3974 <= p3_data_enable ? p2_bit_slice_3974 : p3_bit_slice_3974;
      p3_bit_slice_3975 <= p3_data_enable ? p2_bit_slice_3975 : p3_bit_slice_3975;
      p3_bit_slice_3976 <= p3_data_enable ? p2_bit_slice_3976 : p3_bit_slice_3976;
      p3_bit_slice_3977 <= p3_data_enable ? p2_bit_slice_3977 : p3_bit_slice_3977;
      p3_bit_slice_3978 <= p3_data_enable ? p2_bit_slice_3978 : p3_bit_slice_3978;
      p3_bit_slice_3979 <= p3_data_enable ? p2_bit_slice_3979 : p3_bit_slice_3979;
      p3_bit_slice_3980 <= p3_data_enable ? p2_bit_slice_3980 : p3_bit_slice_3980;
      p3_bit_slice_3981 <= p3_data_enable ? p2_bit_slice_3981 : p3_bit_slice_3981;
      p3_bit_slice_3982 <= p3_data_enable ? p2_bit_slice_3982 : p3_bit_slice_3982;
      p3_bit_slice_3983 <= p3_data_enable ? p2_bit_slice_3983 : p3_bit_slice_3983;
      p3_bit_slice_3984 <= p3_data_enable ? p2_bit_slice_3984 : p3_bit_slice_3984;
      p3_bit_slice_3985 <= p3_data_enable ? p2_bit_slice_3985 : p3_bit_slice_3985;
      p3_bit_slice_3986 <= p3_data_enable ? p2_bit_slice_3986 : p3_bit_slice_3986;
      p3_bit_slice_3987 <= p3_data_enable ? p2_bit_slice_3987 : p3_bit_slice_3987;
      p3_bit_slice_3989 <= p3_data_enable ? p2_bit_slice_3989 : p3_bit_slice_3989;
      p3_bit_slice_3990 <= p3_data_enable ? p2_bit_slice_3990 : p3_bit_slice_3990;
      p3_flag_zero <= p3_data_enable ? flag_zero : p3_flag_zero;
      p3_result_sign <= p3_data_enable ? p2_result_sign : p3_result_sign;
      p3_result_exp <= p3_data_enable ? result_exp : p3_result_exp;
      p4_b_fraction <= p4_data_enable ? p3_b_fraction : p4_b_fraction;
      p4_uge_4116 <= p4_data_enable ? p3_uge_4116 : p4_uge_4116;
      p4_b_fractionivisor__1 <= p4_data_enable ? p3_b_fractionivisor__1 : p4_b_fractionivisor__1;
      p4_uge_4124 <= p4_data_enable ? p3_uge_4124 : p4_uge_4124;
      p4_uge_4195 <= p4_data_enable ? p3_uge_4195 : p4_uge_4195;
      p4_concat_4269 <= p4_data_enable ? concat_4269 : p4_concat_4269;
      p4_uge_4270 <= p4_data_enable ? uge_4270 : p4_uge_4270;
      p4_bit_slice_3971 <= p4_data_enable ? p3_bit_slice_3971 : p4_bit_slice_3971;
      p4_bit_slice_3972 <= p4_data_enable ? p3_bit_slice_3972 : p4_bit_slice_3972;
      p4_bit_slice_3973 <= p4_data_enable ? p3_bit_slice_3973 : p4_bit_slice_3973;
      p4_bit_slice_3974 <= p4_data_enable ? p3_bit_slice_3974 : p4_bit_slice_3974;
      p4_bit_slice_3975 <= p4_data_enable ? p3_bit_slice_3975 : p4_bit_slice_3975;
      p4_bit_slice_3976 <= p4_data_enable ? p3_bit_slice_3976 : p4_bit_slice_3976;
      p4_bit_slice_3977 <= p4_data_enable ? p3_bit_slice_3977 : p4_bit_slice_3977;
      p4_bit_slice_3978 <= p4_data_enable ? p3_bit_slice_3978 : p4_bit_slice_3978;
      p4_bit_slice_3979 <= p4_data_enable ? p3_bit_slice_3979 : p4_bit_slice_3979;
      p4_bit_slice_3980 <= p4_data_enable ? p3_bit_slice_3980 : p4_bit_slice_3980;
      p4_bit_slice_3981 <= p4_data_enable ? p3_bit_slice_3981 : p4_bit_slice_3981;
      p4_bit_slice_3982 <= p4_data_enable ? p3_bit_slice_3982 : p4_bit_slice_3982;
      p4_bit_slice_3983 <= p4_data_enable ? p3_bit_slice_3983 : p4_bit_slice_3983;
      p4_bit_slice_3984 <= p4_data_enable ? p3_bit_slice_3984 : p4_bit_slice_3984;
      p4_bit_slice_3985 <= p4_data_enable ? p3_bit_slice_3985 : p4_bit_slice_3985;
      p4_bit_slice_3986 <= p4_data_enable ? p3_bit_slice_3986 : p4_bit_slice_3986;
      p4_bit_slice_3987 <= p4_data_enable ? p3_bit_slice_3987 : p4_bit_slice_3987;
      p4_bit_slice_3989 <= p4_data_enable ? p3_bit_slice_3989 : p4_bit_slice_3989;
      p4_bit_slice_3990 <= p4_data_enable ? p3_bit_slice_3990 : p4_bit_slice_3990;
      p4_flag_zero <= p4_data_enable ? p3_flag_zero : p4_flag_zero;
      p4_result_sign <= p4_data_enable ? p3_result_sign : p4_result_sign;
      p4_result_exp <= p4_data_enable ? p3_result_exp : p4_result_exp;
      p5_b_fraction <= p5_data_enable ? p4_b_fraction : p5_b_fraction;
      p5_uge_4116 <= p5_data_enable ? p4_uge_4116 : p5_uge_4116;
      p5_b_fractionivisor__1 <= p5_data_enable ? p4_b_fractionivisor__1 : p5_b_fractionivisor__1;
      p5_uge_4124 <= p5_data_enable ? p4_uge_4124 : p5_uge_4124;
      p5_uge_4195 <= p5_data_enable ? p4_uge_4195 : p5_uge_4195;
      p5_uge_4270 <= p5_data_enable ? p4_uge_4270 : p5_uge_4270;
      p5_concat_4335 <= p5_data_enable ? concat_4335 : p5_concat_4335;
      p5_uge_4336 <= p5_data_enable ? uge_4336 : p5_uge_4336;
      p5_bit_slice_3972 <= p5_data_enable ? p4_bit_slice_3972 : p5_bit_slice_3972;
      p5_bit_slice_3973 <= p5_data_enable ? p4_bit_slice_3973 : p5_bit_slice_3973;
      p5_bit_slice_3974 <= p5_data_enable ? p4_bit_slice_3974 : p5_bit_slice_3974;
      p5_bit_slice_3975 <= p5_data_enable ? p4_bit_slice_3975 : p5_bit_slice_3975;
      p5_bit_slice_3976 <= p5_data_enable ? p4_bit_slice_3976 : p5_bit_slice_3976;
      p5_bit_slice_3977 <= p5_data_enable ? p4_bit_slice_3977 : p5_bit_slice_3977;
      p5_bit_slice_3978 <= p5_data_enable ? p4_bit_slice_3978 : p5_bit_slice_3978;
      p5_bit_slice_3979 <= p5_data_enable ? p4_bit_slice_3979 : p5_bit_slice_3979;
      p5_bit_slice_3980 <= p5_data_enable ? p4_bit_slice_3980 : p5_bit_slice_3980;
      p5_bit_slice_3981 <= p5_data_enable ? p4_bit_slice_3981 : p5_bit_slice_3981;
      p5_bit_slice_3982 <= p5_data_enable ? p4_bit_slice_3982 : p5_bit_slice_3982;
      p5_bit_slice_3983 <= p5_data_enable ? p4_bit_slice_3983 : p5_bit_slice_3983;
      p5_bit_slice_3984 <= p5_data_enable ? p4_bit_slice_3984 : p5_bit_slice_3984;
      p5_bit_slice_3985 <= p5_data_enable ? p4_bit_slice_3985 : p5_bit_slice_3985;
      p5_bit_slice_3986 <= p5_data_enable ? p4_bit_slice_3986 : p5_bit_slice_3986;
      p5_bit_slice_3987 <= p5_data_enable ? p4_bit_slice_3987 : p5_bit_slice_3987;
      p5_bit_slice_3989 <= p5_data_enable ? p4_bit_slice_3989 : p5_bit_slice_3989;
      p5_bit_slice_3990 <= p5_data_enable ? p4_bit_slice_3990 : p5_bit_slice_3990;
      p5_flag_zero <= p5_data_enable ? p4_flag_zero : p5_flag_zero;
      p5_result_sign <= p5_data_enable ? p4_result_sign : p5_result_sign;
      p5_result_exp <= p5_data_enable ? p4_result_exp : p5_result_exp;
      p6_b_fraction <= p6_data_enable ? p5_b_fraction : p6_b_fraction;
      p6_uge_4116 <= p6_data_enable ? p5_uge_4116 : p6_uge_4116;
      p6_b_fractionivisor__1 <= p6_data_enable ? p5_b_fractionivisor__1 : p6_b_fractionivisor__1;
      p6_uge_4124 <= p6_data_enable ? p5_uge_4124 : p6_uge_4124;
      p6_uge_4195 <= p6_data_enable ? p5_uge_4195 : p6_uge_4195;
      p6_uge_4270 <= p6_data_enable ? p5_uge_4270 : p6_uge_4270;
      p6_uge_4336 <= p6_data_enable ? p5_uge_4336 : p6_uge_4336;
      p6_concat_4401 <= p6_data_enable ? concat_4401 : p6_concat_4401;
      p6_uge_4402 <= p6_data_enable ? uge_4402 : p6_uge_4402;
      p6_bit_slice_3973 <= p6_data_enable ? p5_bit_slice_3973 : p6_bit_slice_3973;
      p6_bit_slice_3974 <= p6_data_enable ? p5_bit_slice_3974 : p6_bit_slice_3974;
      p6_bit_slice_3975 <= p6_data_enable ? p5_bit_slice_3975 : p6_bit_slice_3975;
      p6_bit_slice_3976 <= p6_data_enable ? p5_bit_slice_3976 : p6_bit_slice_3976;
      p6_bit_slice_3977 <= p6_data_enable ? p5_bit_slice_3977 : p6_bit_slice_3977;
      p6_bit_slice_3978 <= p6_data_enable ? p5_bit_slice_3978 : p6_bit_slice_3978;
      p6_bit_slice_3979 <= p6_data_enable ? p5_bit_slice_3979 : p6_bit_slice_3979;
      p6_bit_slice_3980 <= p6_data_enable ? p5_bit_slice_3980 : p6_bit_slice_3980;
      p6_bit_slice_3981 <= p6_data_enable ? p5_bit_slice_3981 : p6_bit_slice_3981;
      p6_bit_slice_3982 <= p6_data_enable ? p5_bit_slice_3982 : p6_bit_slice_3982;
      p6_bit_slice_3983 <= p6_data_enable ? p5_bit_slice_3983 : p6_bit_slice_3983;
      p6_bit_slice_3984 <= p6_data_enable ? p5_bit_slice_3984 : p6_bit_slice_3984;
      p6_bit_slice_3985 <= p6_data_enable ? p5_bit_slice_3985 : p6_bit_slice_3985;
      p6_bit_slice_3986 <= p6_data_enable ? p5_bit_slice_3986 : p6_bit_slice_3986;
      p6_bit_slice_3987 <= p6_data_enable ? p5_bit_slice_3987 : p6_bit_slice_3987;
      p6_bit_slice_3989 <= p6_data_enable ? p5_bit_slice_3989 : p6_bit_slice_3989;
      p6_bit_slice_3990 <= p6_data_enable ? p5_bit_slice_3990 : p6_bit_slice_3990;
      p6_flag_zero <= p6_data_enable ? p5_flag_zero : p6_flag_zero;
      p6_result_sign <= p6_data_enable ? p5_result_sign : p6_result_sign;
      p6_result_exp <= p6_data_enable ? p5_result_exp : p6_result_exp;
      p7_b_fraction <= p7_data_enable ? p6_b_fraction : p7_b_fraction;
      p7_uge_4116 <= p7_data_enable ? p6_uge_4116 : p7_uge_4116;
      p7_b_fractionivisor__1 <= p7_data_enable ? p6_b_fractionivisor__1 : p7_b_fractionivisor__1;
      p7_uge_4124 <= p7_data_enable ? p6_uge_4124 : p7_uge_4124;
      p7_uge_4195 <= p7_data_enable ? p6_uge_4195 : p7_uge_4195;
      p7_uge_4270 <= p7_data_enable ? p6_uge_4270 : p7_uge_4270;
      p7_uge_4336 <= p7_data_enable ? p6_uge_4336 : p7_uge_4336;
      p7_uge_4402 <= p7_data_enable ? p6_uge_4402 : p7_uge_4402;
      p7_concat_4467 <= p7_data_enable ? concat_4467 : p7_concat_4467;
      p7_uge_4468 <= p7_data_enable ? uge_4468 : p7_uge_4468;
      p7_bit_slice_3974 <= p7_data_enable ? p6_bit_slice_3974 : p7_bit_slice_3974;
      p7_bit_slice_3975 <= p7_data_enable ? p6_bit_slice_3975 : p7_bit_slice_3975;
      p7_bit_slice_3976 <= p7_data_enable ? p6_bit_slice_3976 : p7_bit_slice_3976;
      p7_bit_slice_3977 <= p7_data_enable ? p6_bit_slice_3977 : p7_bit_slice_3977;
      p7_bit_slice_3978 <= p7_data_enable ? p6_bit_slice_3978 : p7_bit_slice_3978;
      p7_bit_slice_3979 <= p7_data_enable ? p6_bit_slice_3979 : p7_bit_slice_3979;
      p7_bit_slice_3980 <= p7_data_enable ? p6_bit_slice_3980 : p7_bit_slice_3980;
      p7_bit_slice_3981 <= p7_data_enable ? p6_bit_slice_3981 : p7_bit_slice_3981;
      p7_bit_slice_3982 <= p7_data_enable ? p6_bit_slice_3982 : p7_bit_slice_3982;
      p7_bit_slice_3983 <= p7_data_enable ? p6_bit_slice_3983 : p7_bit_slice_3983;
      p7_bit_slice_3984 <= p7_data_enable ? p6_bit_slice_3984 : p7_bit_slice_3984;
      p7_bit_slice_3985 <= p7_data_enable ? p6_bit_slice_3985 : p7_bit_slice_3985;
      p7_bit_slice_3986 <= p7_data_enable ? p6_bit_slice_3986 : p7_bit_slice_3986;
      p7_bit_slice_3987 <= p7_data_enable ? p6_bit_slice_3987 : p7_bit_slice_3987;
      p7_bit_slice_3989 <= p7_data_enable ? p6_bit_slice_3989 : p7_bit_slice_3989;
      p7_bit_slice_3990 <= p7_data_enable ? p6_bit_slice_3990 : p7_bit_slice_3990;
      p7_flag_zero <= p7_data_enable ? p6_flag_zero : p7_flag_zero;
      p7_result_sign <= p7_data_enable ? p6_result_sign : p7_result_sign;
      p7_result_exp <= p7_data_enable ? p6_result_exp : p7_result_exp;
      p8_b_fraction <= p8_data_enable ? p7_b_fraction : p8_b_fraction;
      p8_uge_4116 <= p8_data_enable ? p7_uge_4116 : p8_uge_4116;
      p8_b_fractionivisor__1 <= p8_data_enable ? p7_b_fractionivisor__1 : p8_b_fractionivisor__1;
      p8_uge_4124 <= p8_data_enable ? p7_uge_4124 : p8_uge_4124;
      p8_uge_4195 <= p8_data_enable ? p7_uge_4195 : p8_uge_4195;
      p8_uge_4270 <= p8_data_enable ? p7_uge_4270 : p8_uge_4270;
      p8_uge_4336 <= p8_data_enable ? p7_uge_4336 : p8_uge_4336;
      p8_uge_4402 <= p8_data_enable ? p7_uge_4402 : p8_uge_4402;
      p8_uge_4468 <= p8_data_enable ? p7_uge_4468 : p8_uge_4468;
      p8_concat_4533 <= p8_data_enable ? concat_4533 : p8_concat_4533;
      p8_uge_4534 <= p8_data_enable ? uge_4534 : p8_uge_4534;
      p8_bit_slice_3975 <= p8_data_enable ? p7_bit_slice_3975 : p8_bit_slice_3975;
      p8_bit_slice_3976 <= p8_data_enable ? p7_bit_slice_3976 : p8_bit_slice_3976;
      p8_bit_slice_3977 <= p8_data_enable ? p7_bit_slice_3977 : p8_bit_slice_3977;
      p8_bit_slice_3978 <= p8_data_enable ? p7_bit_slice_3978 : p8_bit_slice_3978;
      p8_bit_slice_3979 <= p8_data_enable ? p7_bit_slice_3979 : p8_bit_slice_3979;
      p8_bit_slice_3980 <= p8_data_enable ? p7_bit_slice_3980 : p8_bit_slice_3980;
      p8_bit_slice_3981 <= p8_data_enable ? p7_bit_slice_3981 : p8_bit_slice_3981;
      p8_bit_slice_3982 <= p8_data_enable ? p7_bit_slice_3982 : p8_bit_slice_3982;
      p8_bit_slice_3983 <= p8_data_enable ? p7_bit_slice_3983 : p8_bit_slice_3983;
      p8_bit_slice_3984 <= p8_data_enable ? p7_bit_slice_3984 : p8_bit_slice_3984;
      p8_bit_slice_3985 <= p8_data_enable ? p7_bit_slice_3985 : p8_bit_slice_3985;
      p8_bit_slice_3986 <= p8_data_enable ? p7_bit_slice_3986 : p8_bit_slice_3986;
      p8_bit_slice_3987 <= p8_data_enable ? p7_bit_slice_3987 : p8_bit_slice_3987;
      p8_bit_slice_3989 <= p8_data_enable ? p7_bit_slice_3989 : p8_bit_slice_3989;
      p8_bit_slice_3990 <= p8_data_enable ? p7_bit_slice_3990 : p8_bit_slice_3990;
      p8_flag_zero <= p8_data_enable ? p7_flag_zero : p8_flag_zero;
      p8_result_sign <= p8_data_enable ? p7_result_sign : p8_result_sign;
      p8_result_exp <= p8_data_enable ? p7_result_exp : p8_result_exp;
      p9_b_fraction <= p9_data_enable ? p8_b_fraction : p9_b_fraction;
      p9_uge_4116 <= p9_data_enable ? p8_uge_4116 : p9_uge_4116;
      p9_b_fractionivisor__1 <= p9_data_enable ? p8_b_fractionivisor__1 : p9_b_fractionivisor__1;
      p9_uge_4124 <= p9_data_enable ? p8_uge_4124 : p9_uge_4124;
      p9_uge_4195 <= p9_data_enable ? p8_uge_4195 : p9_uge_4195;
      p9_uge_4270 <= p9_data_enable ? p8_uge_4270 : p9_uge_4270;
      p9_uge_4336 <= p9_data_enable ? p8_uge_4336 : p9_uge_4336;
      p9_uge_4402 <= p9_data_enable ? p8_uge_4402 : p9_uge_4402;
      p9_uge_4468 <= p9_data_enable ? p8_uge_4468 : p9_uge_4468;
      p9_uge_4534 <= p9_data_enable ? p8_uge_4534 : p9_uge_4534;
      p9_concat_4599 <= p9_data_enable ? concat_4599 : p9_concat_4599;
      p9_uge_4600 <= p9_data_enable ? uge_4600 : p9_uge_4600;
      p9_bit_slice_3976 <= p9_data_enable ? p8_bit_slice_3976 : p9_bit_slice_3976;
      p9_bit_slice_3977 <= p9_data_enable ? p8_bit_slice_3977 : p9_bit_slice_3977;
      p9_bit_slice_3978 <= p9_data_enable ? p8_bit_slice_3978 : p9_bit_slice_3978;
      p9_bit_slice_3979 <= p9_data_enable ? p8_bit_slice_3979 : p9_bit_slice_3979;
      p9_bit_slice_3980 <= p9_data_enable ? p8_bit_slice_3980 : p9_bit_slice_3980;
      p9_bit_slice_3981 <= p9_data_enable ? p8_bit_slice_3981 : p9_bit_slice_3981;
      p9_bit_slice_3982 <= p9_data_enable ? p8_bit_slice_3982 : p9_bit_slice_3982;
      p9_bit_slice_3983 <= p9_data_enable ? p8_bit_slice_3983 : p9_bit_slice_3983;
      p9_bit_slice_3984 <= p9_data_enable ? p8_bit_slice_3984 : p9_bit_slice_3984;
      p9_bit_slice_3985 <= p9_data_enable ? p8_bit_slice_3985 : p9_bit_slice_3985;
      p9_bit_slice_3986 <= p9_data_enable ? p8_bit_slice_3986 : p9_bit_slice_3986;
      p9_bit_slice_3987 <= p9_data_enable ? p8_bit_slice_3987 : p9_bit_slice_3987;
      p9_bit_slice_3989 <= p9_data_enable ? p8_bit_slice_3989 : p9_bit_slice_3989;
      p9_bit_slice_3990 <= p9_data_enable ? p8_bit_slice_3990 : p9_bit_slice_3990;
      p9_flag_zero <= p9_data_enable ? p8_flag_zero : p9_flag_zero;
      p9_result_sign <= p9_data_enable ? p8_result_sign : p9_result_sign;
      p9_result_exp <= p9_data_enable ? p8_result_exp : p9_result_exp;
      p10_b_fraction <= p10_data_enable ? p9_b_fraction : p10_b_fraction;
      p10_uge_4116 <= p10_data_enable ? p9_uge_4116 : p10_uge_4116;
      p10_b_fractionivisor__1 <= p10_data_enable ? p9_b_fractionivisor__1 : p10_b_fractionivisor__1;
      p10_uge_4124 <= p10_data_enable ? p9_uge_4124 : p10_uge_4124;
      p10_uge_4195 <= p10_data_enable ? p9_uge_4195 : p10_uge_4195;
      p10_uge_4270 <= p10_data_enable ? p9_uge_4270 : p10_uge_4270;
      p10_uge_4336 <= p10_data_enable ? p9_uge_4336 : p10_uge_4336;
      p10_uge_4402 <= p10_data_enable ? p9_uge_4402 : p10_uge_4402;
      p10_uge_4468 <= p10_data_enable ? p9_uge_4468 : p10_uge_4468;
      p10_uge_4534 <= p10_data_enable ? p9_uge_4534 : p10_uge_4534;
      p10_uge_4600 <= p10_data_enable ? p9_uge_4600 : p10_uge_4600;
      p10_concat_4665 <= p10_data_enable ? concat_4665 : p10_concat_4665;
      p10_uge_4666 <= p10_data_enable ? uge_4666 : p10_uge_4666;
      p10_bit_slice_3977 <= p10_data_enable ? p9_bit_slice_3977 : p10_bit_slice_3977;
      p10_bit_slice_3978 <= p10_data_enable ? p9_bit_slice_3978 : p10_bit_slice_3978;
      p10_bit_slice_3979 <= p10_data_enable ? p9_bit_slice_3979 : p10_bit_slice_3979;
      p10_bit_slice_3980 <= p10_data_enable ? p9_bit_slice_3980 : p10_bit_slice_3980;
      p10_bit_slice_3981 <= p10_data_enable ? p9_bit_slice_3981 : p10_bit_slice_3981;
      p10_bit_slice_3982 <= p10_data_enable ? p9_bit_slice_3982 : p10_bit_slice_3982;
      p10_bit_slice_3983 <= p10_data_enable ? p9_bit_slice_3983 : p10_bit_slice_3983;
      p10_bit_slice_3984 <= p10_data_enable ? p9_bit_slice_3984 : p10_bit_slice_3984;
      p10_bit_slice_3985 <= p10_data_enable ? p9_bit_slice_3985 : p10_bit_slice_3985;
      p10_bit_slice_3986 <= p10_data_enable ? p9_bit_slice_3986 : p10_bit_slice_3986;
      p10_bit_slice_3987 <= p10_data_enable ? p9_bit_slice_3987 : p10_bit_slice_3987;
      p10_bit_slice_3989 <= p10_data_enable ? p9_bit_slice_3989 : p10_bit_slice_3989;
      p10_bit_slice_3990 <= p10_data_enable ? p9_bit_slice_3990 : p10_bit_slice_3990;
      p10_flag_zero <= p10_data_enable ? p9_flag_zero : p10_flag_zero;
      p10_result_sign <= p10_data_enable ? p9_result_sign : p10_result_sign;
      p10_result_exp <= p10_data_enable ? p9_result_exp : p10_result_exp;
      p11_b_fraction <= p11_data_enable ? p10_b_fraction : p11_b_fraction;
      p11_uge_4116 <= p11_data_enable ? p10_uge_4116 : p11_uge_4116;
      p11_b_fractionivisor__1 <= p11_data_enable ? p10_b_fractionivisor__1 : p11_b_fractionivisor__1;
      p11_uge_4124 <= p11_data_enable ? p10_uge_4124 : p11_uge_4124;
      p11_uge_4195 <= p11_data_enable ? p10_uge_4195 : p11_uge_4195;
      p11_uge_4270 <= p11_data_enable ? p10_uge_4270 : p11_uge_4270;
      p11_uge_4336 <= p11_data_enable ? p10_uge_4336 : p11_uge_4336;
      p11_uge_4402 <= p11_data_enable ? p10_uge_4402 : p11_uge_4402;
      p11_uge_4468 <= p11_data_enable ? p10_uge_4468 : p11_uge_4468;
      p11_uge_4534 <= p11_data_enable ? p10_uge_4534 : p11_uge_4534;
      p11_uge_4600 <= p11_data_enable ? p10_uge_4600 : p11_uge_4600;
      p11_uge_4666 <= p11_data_enable ? p10_uge_4666 : p11_uge_4666;
      p11_concat_4731 <= p11_data_enable ? concat_4731 : p11_concat_4731;
      p11_uge_4732 <= p11_data_enable ? uge_4732 : p11_uge_4732;
      p11_bit_slice_3978 <= p11_data_enable ? p10_bit_slice_3978 : p11_bit_slice_3978;
      p11_bit_slice_3979 <= p11_data_enable ? p10_bit_slice_3979 : p11_bit_slice_3979;
      p11_bit_slice_3980 <= p11_data_enable ? p10_bit_slice_3980 : p11_bit_slice_3980;
      p11_bit_slice_3981 <= p11_data_enable ? p10_bit_slice_3981 : p11_bit_slice_3981;
      p11_bit_slice_3982 <= p11_data_enable ? p10_bit_slice_3982 : p11_bit_slice_3982;
      p11_bit_slice_3983 <= p11_data_enable ? p10_bit_slice_3983 : p11_bit_slice_3983;
      p11_bit_slice_3984 <= p11_data_enable ? p10_bit_slice_3984 : p11_bit_slice_3984;
      p11_bit_slice_3985 <= p11_data_enable ? p10_bit_slice_3985 : p11_bit_slice_3985;
      p11_bit_slice_3986 <= p11_data_enable ? p10_bit_slice_3986 : p11_bit_slice_3986;
      p11_bit_slice_3987 <= p11_data_enable ? p10_bit_slice_3987 : p11_bit_slice_3987;
      p11_bit_slice_3989 <= p11_data_enable ? p10_bit_slice_3989 : p11_bit_slice_3989;
      p11_bit_slice_3990 <= p11_data_enable ? p10_bit_slice_3990 : p11_bit_slice_3990;
      p11_flag_zero <= p11_data_enable ? p10_flag_zero : p11_flag_zero;
      p11_result_sign <= p11_data_enable ? p10_result_sign : p11_result_sign;
      p11_result_exp <= p11_data_enable ? p10_result_exp : p11_result_exp;
      p12_b_fraction <= p12_data_enable ? p11_b_fraction : p12_b_fraction;
      p12_uge_4116 <= p12_data_enable ? p11_uge_4116 : p12_uge_4116;
      p12_b_fractionivisor__1 <= p12_data_enable ? p11_b_fractionivisor__1 : p12_b_fractionivisor__1;
      p12_uge_4124 <= p12_data_enable ? p11_uge_4124 : p12_uge_4124;
      p12_uge_4195 <= p12_data_enable ? p11_uge_4195 : p12_uge_4195;
      p12_uge_4270 <= p12_data_enable ? p11_uge_4270 : p12_uge_4270;
      p12_uge_4336 <= p12_data_enable ? p11_uge_4336 : p12_uge_4336;
      p12_uge_4402 <= p12_data_enable ? p11_uge_4402 : p12_uge_4402;
      p12_uge_4468 <= p12_data_enable ? p11_uge_4468 : p12_uge_4468;
      p12_uge_4534 <= p12_data_enable ? p11_uge_4534 : p12_uge_4534;
      p12_uge_4600 <= p12_data_enable ? p11_uge_4600 : p12_uge_4600;
      p12_uge_4666 <= p12_data_enable ? p11_uge_4666 : p12_uge_4666;
      p12_uge_4732 <= p12_data_enable ? p11_uge_4732 : p12_uge_4732;
      p12_concat_4797 <= p12_data_enable ? concat_4797 : p12_concat_4797;
      p12_uge_4798 <= p12_data_enable ? uge_4798 : p12_uge_4798;
      p12_bit_slice_3979 <= p12_data_enable ? p11_bit_slice_3979 : p12_bit_slice_3979;
      p12_bit_slice_3980 <= p12_data_enable ? p11_bit_slice_3980 : p12_bit_slice_3980;
      p12_bit_slice_3981 <= p12_data_enable ? p11_bit_slice_3981 : p12_bit_slice_3981;
      p12_bit_slice_3982 <= p12_data_enable ? p11_bit_slice_3982 : p12_bit_slice_3982;
      p12_bit_slice_3983 <= p12_data_enable ? p11_bit_slice_3983 : p12_bit_slice_3983;
      p12_bit_slice_3984 <= p12_data_enable ? p11_bit_slice_3984 : p12_bit_slice_3984;
      p12_bit_slice_3985 <= p12_data_enable ? p11_bit_slice_3985 : p12_bit_slice_3985;
      p12_bit_slice_3986 <= p12_data_enable ? p11_bit_slice_3986 : p12_bit_slice_3986;
      p12_bit_slice_3987 <= p12_data_enable ? p11_bit_slice_3987 : p12_bit_slice_3987;
      p12_bit_slice_3989 <= p12_data_enable ? p11_bit_slice_3989 : p12_bit_slice_3989;
      p12_bit_slice_3990 <= p12_data_enable ? p11_bit_slice_3990 : p12_bit_slice_3990;
      p12_flag_zero <= p12_data_enable ? p11_flag_zero : p12_flag_zero;
      p12_result_sign <= p12_data_enable ? p11_result_sign : p12_result_sign;
      p12_result_exp <= p12_data_enable ? p11_result_exp : p12_result_exp;
      p13_b_fraction <= p13_data_enable ? p12_b_fraction : p13_b_fraction;
      p13_uge_4116 <= p13_data_enable ? p12_uge_4116 : p13_uge_4116;
      p13_b_fractionivisor__1 <= p13_data_enable ? p12_b_fractionivisor__1 : p13_b_fractionivisor__1;
      p13_uge_4124 <= p13_data_enable ? p12_uge_4124 : p13_uge_4124;
      p13_uge_4195 <= p13_data_enable ? p12_uge_4195 : p13_uge_4195;
      p13_uge_4270 <= p13_data_enable ? p12_uge_4270 : p13_uge_4270;
      p13_uge_4336 <= p13_data_enable ? p12_uge_4336 : p13_uge_4336;
      p13_uge_4402 <= p13_data_enable ? p12_uge_4402 : p13_uge_4402;
      p13_uge_4468 <= p13_data_enable ? p12_uge_4468 : p13_uge_4468;
      p13_uge_4534 <= p13_data_enable ? p12_uge_4534 : p13_uge_4534;
      p13_uge_4600 <= p13_data_enable ? p12_uge_4600 : p13_uge_4600;
      p13_uge_4666 <= p13_data_enable ? p12_uge_4666 : p13_uge_4666;
      p13_uge_4732 <= p13_data_enable ? p12_uge_4732 : p13_uge_4732;
      p13_uge_4798 <= p13_data_enable ? p12_uge_4798 : p13_uge_4798;
      p13_concat_4863 <= p13_data_enable ? concat_4863 : p13_concat_4863;
      p13_uge_4864 <= p13_data_enable ? uge_4864 : p13_uge_4864;
      p13_bit_slice_3980 <= p13_data_enable ? p12_bit_slice_3980 : p13_bit_slice_3980;
      p13_bit_slice_3981 <= p13_data_enable ? p12_bit_slice_3981 : p13_bit_slice_3981;
      p13_bit_slice_3982 <= p13_data_enable ? p12_bit_slice_3982 : p13_bit_slice_3982;
      p13_bit_slice_3983 <= p13_data_enable ? p12_bit_slice_3983 : p13_bit_slice_3983;
      p13_bit_slice_3984 <= p13_data_enable ? p12_bit_slice_3984 : p13_bit_slice_3984;
      p13_bit_slice_3985 <= p13_data_enable ? p12_bit_slice_3985 : p13_bit_slice_3985;
      p13_bit_slice_3986 <= p13_data_enable ? p12_bit_slice_3986 : p13_bit_slice_3986;
      p13_bit_slice_3987 <= p13_data_enable ? p12_bit_slice_3987 : p13_bit_slice_3987;
      p13_bit_slice_3989 <= p13_data_enable ? p12_bit_slice_3989 : p13_bit_slice_3989;
      p13_bit_slice_3990 <= p13_data_enable ? p12_bit_slice_3990 : p13_bit_slice_3990;
      p13_flag_zero <= p13_data_enable ? p12_flag_zero : p13_flag_zero;
      p13_result_sign <= p13_data_enable ? p12_result_sign : p13_result_sign;
      p13_result_exp <= p13_data_enable ? p12_result_exp : p13_result_exp;
      p14_b_fraction <= p14_data_enable ? p13_b_fraction : p14_b_fraction;
      p14_uge_4116 <= p14_data_enable ? p13_uge_4116 : p14_uge_4116;
      p14_b_fractionivisor__1 <= p14_data_enable ? p13_b_fractionivisor__1 : p14_b_fractionivisor__1;
      p14_uge_4124 <= p14_data_enable ? p13_uge_4124 : p14_uge_4124;
      p14_uge_4195 <= p14_data_enable ? p13_uge_4195 : p14_uge_4195;
      p14_uge_4270 <= p14_data_enable ? p13_uge_4270 : p14_uge_4270;
      p14_uge_4336 <= p14_data_enable ? p13_uge_4336 : p14_uge_4336;
      p14_uge_4402 <= p14_data_enable ? p13_uge_4402 : p14_uge_4402;
      p14_uge_4468 <= p14_data_enable ? p13_uge_4468 : p14_uge_4468;
      p14_uge_4534 <= p14_data_enable ? p13_uge_4534 : p14_uge_4534;
      p14_uge_4600 <= p14_data_enable ? p13_uge_4600 : p14_uge_4600;
      p14_uge_4666 <= p14_data_enable ? p13_uge_4666 : p14_uge_4666;
      p14_uge_4732 <= p14_data_enable ? p13_uge_4732 : p14_uge_4732;
      p14_uge_4798 <= p14_data_enable ? p13_uge_4798 : p14_uge_4798;
      p14_uge_4864 <= p14_data_enable ? p13_uge_4864 : p14_uge_4864;
      p14_concat_4929 <= p14_data_enable ? concat_4929 : p14_concat_4929;
      p14_uge_4930 <= p14_data_enable ? uge_4930 : p14_uge_4930;
      p14_bit_slice_3981 <= p14_data_enable ? p13_bit_slice_3981 : p14_bit_slice_3981;
      p14_bit_slice_3982 <= p14_data_enable ? p13_bit_slice_3982 : p14_bit_slice_3982;
      p14_bit_slice_3983 <= p14_data_enable ? p13_bit_slice_3983 : p14_bit_slice_3983;
      p14_bit_slice_3984 <= p14_data_enable ? p13_bit_slice_3984 : p14_bit_slice_3984;
      p14_bit_slice_3985 <= p14_data_enable ? p13_bit_slice_3985 : p14_bit_slice_3985;
      p14_bit_slice_3986 <= p14_data_enable ? p13_bit_slice_3986 : p14_bit_slice_3986;
      p14_bit_slice_3987 <= p14_data_enable ? p13_bit_slice_3987 : p14_bit_slice_3987;
      p14_bit_slice_3989 <= p14_data_enable ? p13_bit_slice_3989 : p14_bit_slice_3989;
      p14_bit_slice_3990 <= p14_data_enable ? p13_bit_slice_3990 : p14_bit_slice_3990;
      p14_flag_zero <= p14_data_enable ? p13_flag_zero : p14_flag_zero;
      p14_result_sign <= p14_data_enable ? p13_result_sign : p14_result_sign;
      p14_result_exp <= p14_data_enable ? p13_result_exp : p14_result_exp;
      p15_b_fraction <= p15_data_enable ? p14_b_fraction : p15_b_fraction;
      p15_uge_4116 <= p15_data_enable ? p14_uge_4116 : p15_uge_4116;
      p15_b_fractionivisor__1 <= p15_data_enable ? p14_b_fractionivisor__1 : p15_b_fractionivisor__1;
      p15_uge_4124 <= p15_data_enable ? p14_uge_4124 : p15_uge_4124;
      p15_uge_4195 <= p15_data_enable ? p14_uge_4195 : p15_uge_4195;
      p15_uge_4270 <= p15_data_enable ? p14_uge_4270 : p15_uge_4270;
      p15_uge_4336 <= p15_data_enable ? p14_uge_4336 : p15_uge_4336;
      p15_uge_4402 <= p15_data_enable ? p14_uge_4402 : p15_uge_4402;
      p15_uge_4468 <= p15_data_enable ? p14_uge_4468 : p15_uge_4468;
      p15_uge_4534 <= p15_data_enable ? p14_uge_4534 : p15_uge_4534;
      p15_uge_4600 <= p15_data_enable ? p14_uge_4600 : p15_uge_4600;
      p15_uge_4666 <= p15_data_enable ? p14_uge_4666 : p15_uge_4666;
      p15_uge_4732 <= p15_data_enable ? p14_uge_4732 : p15_uge_4732;
      p15_uge_4798 <= p15_data_enable ? p14_uge_4798 : p15_uge_4798;
      p15_uge_4864 <= p15_data_enable ? p14_uge_4864 : p15_uge_4864;
      p15_uge_4930 <= p15_data_enable ? p14_uge_4930 : p15_uge_4930;
      p15_concat_4995 <= p15_data_enable ? concat_4995 : p15_concat_4995;
      p15_uge_4996 <= p15_data_enable ? uge_4996 : p15_uge_4996;
      p15_bit_slice_3982 <= p15_data_enable ? p14_bit_slice_3982 : p15_bit_slice_3982;
      p15_bit_slice_3983 <= p15_data_enable ? p14_bit_slice_3983 : p15_bit_slice_3983;
      p15_bit_slice_3984 <= p15_data_enable ? p14_bit_slice_3984 : p15_bit_slice_3984;
      p15_bit_slice_3985 <= p15_data_enable ? p14_bit_slice_3985 : p15_bit_slice_3985;
      p15_bit_slice_3986 <= p15_data_enable ? p14_bit_slice_3986 : p15_bit_slice_3986;
      p15_bit_slice_3987 <= p15_data_enable ? p14_bit_slice_3987 : p15_bit_slice_3987;
      p15_bit_slice_3989 <= p15_data_enable ? p14_bit_slice_3989 : p15_bit_slice_3989;
      p15_bit_slice_3990 <= p15_data_enable ? p14_bit_slice_3990 : p15_bit_slice_3990;
      p15_flag_zero <= p15_data_enable ? p14_flag_zero : p15_flag_zero;
      p15_result_sign <= p15_data_enable ? p14_result_sign : p15_result_sign;
      p15_result_exp <= p15_data_enable ? p14_result_exp : p15_result_exp;
      p16_b_fraction <= p16_data_enable ? p15_b_fraction : p16_b_fraction;
      p16_uge_4116 <= p16_data_enable ? p15_uge_4116 : p16_uge_4116;
      p16_b_fractionivisor__1 <= p16_data_enable ? p15_b_fractionivisor__1 : p16_b_fractionivisor__1;
      p16_uge_4124 <= p16_data_enable ? p15_uge_4124 : p16_uge_4124;
      p16_uge_4195 <= p16_data_enable ? p15_uge_4195 : p16_uge_4195;
      p16_uge_4270 <= p16_data_enable ? p15_uge_4270 : p16_uge_4270;
      p16_uge_4336 <= p16_data_enable ? p15_uge_4336 : p16_uge_4336;
      p16_uge_4402 <= p16_data_enable ? p15_uge_4402 : p16_uge_4402;
      p16_uge_4468 <= p16_data_enable ? p15_uge_4468 : p16_uge_4468;
      p16_uge_4534 <= p16_data_enable ? p15_uge_4534 : p16_uge_4534;
      p16_uge_4600 <= p16_data_enable ? p15_uge_4600 : p16_uge_4600;
      p16_uge_4666 <= p16_data_enable ? p15_uge_4666 : p16_uge_4666;
      p16_uge_4732 <= p16_data_enable ? p15_uge_4732 : p16_uge_4732;
      p16_uge_4798 <= p16_data_enable ? p15_uge_4798 : p16_uge_4798;
      p16_uge_4864 <= p16_data_enable ? p15_uge_4864 : p16_uge_4864;
      p16_uge_4930 <= p16_data_enable ? p15_uge_4930 : p16_uge_4930;
      p16_uge_4996 <= p16_data_enable ? p15_uge_4996 : p16_uge_4996;
      p16_concat_5061 <= p16_data_enable ? concat_5061 : p16_concat_5061;
      p16_uge_5062 <= p16_data_enable ? uge_5062 : p16_uge_5062;
      p16_bit_slice_3983 <= p16_data_enable ? p15_bit_slice_3983 : p16_bit_slice_3983;
      p16_bit_slice_3984 <= p16_data_enable ? p15_bit_slice_3984 : p16_bit_slice_3984;
      p16_bit_slice_3985 <= p16_data_enable ? p15_bit_slice_3985 : p16_bit_slice_3985;
      p16_bit_slice_3986 <= p16_data_enable ? p15_bit_slice_3986 : p16_bit_slice_3986;
      p16_bit_slice_3987 <= p16_data_enable ? p15_bit_slice_3987 : p16_bit_slice_3987;
      p16_bit_slice_3989 <= p16_data_enable ? p15_bit_slice_3989 : p16_bit_slice_3989;
      p16_bit_slice_3990 <= p16_data_enable ? p15_bit_slice_3990 : p16_bit_slice_3990;
      p16_flag_zero <= p16_data_enable ? p15_flag_zero : p16_flag_zero;
      p16_result_sign <= p16_data_enable ? p15_result_sign : p16_result_sign;
      p16_result_exp <= p16_data_enable ? p15_result_exp : p16_result_exp;
      p17_b_fraction <= p17_data_enable ? p16_b_fraction : p17_b_fraction;
      p17_uge_4116 <= p17_data_enable ? p16_uge_4116 : p17_uge_4116;
      p17_b_fractionivisor__1 <= p17_data_enable ? p16_b_fractionivisor__1 : p17_b_fractionivisor__1;
      p17_uge_4124 <= p17_data_enable ? p16_uge_4124 : p17_uge_4124;
      p17_uge_4195 <= p17_data_enable ? p16_uge_4195 : p17_uge_4195;
      p17_uge_4270 <= p17_data_enable ? p16_uge_4270 : p17_uge_4270;
      p17_uge_4336 <= p17_data_enable ? p16_uge_4336 : p17_uge_4336;
      p17_uge_4402 <= p17_data_enable ? p16_uge_4402 : p17_uge_4402;
      p17_uge_4468 <= p17_data_enable ? p16_uge_4468 : p17_uge_4468;
      p17_uge_4534 <= p17_data_enable ? p16_uge_4534 : p17_uge_4534;
      p17_uge_4600 <= p17_data_enable ? p16_uge_4600 : p17_uge_4600;
      p17_uge_4666 <= p17_data_enable ? p16_uge_4666 : p17_uge_4666;
      p17_uge_4732 <= p17_data_enable ? p16_uge_4732 : p17_uge_4732;
      p17_uge_4798 <= p17_data_enable ? p16_uge_4798 : p17_uge_4798;
      p17_uge_4864 <= p17_data_enable ? p16_uge_4864 : p17_uge_4864;
      p17_uge_4930 <= p17_data_enable ? p16_uge_4930 : p17_uge_4930;
      p17_uge_4996 <= p17_data_enable ? p16_uge_4996 : p17_uge_4996;
      p17_uge_5062 <= p17_data_enable ? p16_uge_5062 : p17_uge_5062;
      p17_concat_5127 <= p17_data_enable ? concat_5127 : p17_concat_5127;
      p17_uge_5128 <= p17_data_enable ? uge_5128 : p17_uge_5128;
      p17_bit_slice_3984 <= p17_data_enable ? p16_bit_slice_3984 : p17_bit_slice_3984;
      p17_bit_slice_3985 <= p17_data_enable ? p16_bit_slice_3985 : p17_bit_slice_3985;
      p17_bit_slice_3986 <= p17_data_enable ? p16_bit_slice_3986 : p17_bit_slice_3986;
      p17_bit_slice_3987 <= p17_data_enable ? p16_bit_slice_3987 : p17_bit_slice_3987;
      p17_bit_slice_3989 <= p17_data_enable ? p16_bit_slice_3989 : p17_bit_slice_3989;
      p17_bit_slice_3990 <= p17_data_enable ? p16_bit_slice_3990 : p17_bit_slice_3990;
      p17_flag_zero <= p17_data_enable ? p16_flag_zero : p17_flag_zero;
      p17_result_sign <= p17_data_enable ? p16_result_sign : p17_result_sign;
      p17_result_exp <= p17_data_enable ? p16_result_exp : p17_result_exp;
      p18_b_fraction <= p18_data_enable ? p17_b_fraction : p18_b_fraction;
      p18_uge_4116 <= p18_data_enable ? p17_uge_4116 : p18_uge_4116;
      p18_b_fractionivisor__1 <= p18_data_enable ? p17_b_fractionivisor__1 : p18_b_fractionivisor__1;
      p18_uge_4124 <= p18_data_enable ? p17_uge_4124 : p18_uge_4124;
      p18_uge_4195 <= p18_data_enable ? p17_uge_4195 : p18_uge_4195;
      p18_uge_4270 <= p18_data_enable ? p17_uge_4270 : p18_uge_4270;
      p18_uge_4336 <= p18_data_enable ? p17_uge_4336 : p18_uge_4336;
      p18_uge_4402 <= p18_data_enable ? p17_uge_4402 : p18_uge_4402;
      p18_uge_4468 <= p18_data_enable ? p17_uge_4468 : p18_uge_4468;
      p18_uge_4534 <= p18_data_enable ? p17_uge_4534 : p18_uge_4534;
      p18_uge_4600 <= p18_data_enable ? p17_uge_4600 : p18_uge_4600;
      p18_uge_4666 <= p18_data_enable ? p17_uge_4666 : p18_uge_4666;
      p18_uge_4732 <= p18_data_enable ? p17_uge_4732 : p18_uge_4732;
      p18_uge_4798 <= p18_data_enable ? p17_uge_4798 : p18_uge_4798;
      p18_uge_4864 <= p18_data_enable ? p17_uge_4864 : p18_uge_4864;
      p18_uge_4930 <= p18_data_enable ? p17_uge_4930 : p18_uge_4930;
      p18_uge_4996 <= p18_data_enable ? p17_uge_4996 : p18_uge_4996;
      p18_uge_5062 <= p18_data_enable ? p17_uge_5062 : p18_uge_5062;
      p18_uge_5128 <= p18_data_enable ? p17_uge_5128 : p18_uge_5128;
      p18_concat_5193 <= p18_data_enable ? concat_5193 : p18_concat_5193;
      p18_uge_5194 <= p18_data_enable ? uge_5194 : p18_uge_5194;
      p18_bit_slice_3985 <= p18_data_enable ? p17_bit_slice_3985 : p18_bit_slice_3985;
      p18_bit_slice_3986 <= p18_data_enable ? p17_bit_slice_3986 : p18_bit_slice_3986;
      p18_bit_slice_3987 <= p18_data_enable ? p17_bit_slice_3987 : p18_bit_slice_3987;
      p18_bit_slice_3989 <= p18_data_enable ? p17_bit_slice_3989 : p18_bit_slice_3989;
      p18_bit_slice_3990 <= p18_data_enable ? p17_bit_slice_3990 : p18_bit_slice_3990;
      p18_flag_zero <= p18_data_enable ? p17_flag_zero : p18_flag_zero;
      p18_result_sign <= p18_data_enable ? p17_result_sign : p18_result_sign;
      p18_result_exp <= p18_data_enable ? p17_result_exp : p18_result_exp;
      p19_b_fraction <= p19_data_enable ? p18_b_fraction : p19_b_fraction;
      p19_uge_4116 <= p19_data_enable ? p18_uge_4116 : p19_uge_4116;
      p19_b_fractionivisor__1 <= p19_data_enable ? p18_b_fractionivisor__1 : p19_b_fractionivisor__1;
      p19_uge_4124 <= p19_data_enable ? p18_uge_4124 : p19_uge_4124;
      p19_uge_4195 <= p19_data_enable ? p18_uge_4195 : p19_uge_4195;
      p19_uge_4270 <= p19_data_enable ? p18_uge_4270 : p19_uge_4270;
      p19_uge_4336 <= p19_data_enable ? p18_uge_4336 : p19_uge_4336;
      p19_uge_4402 <= p19_data_enable ? p18_uge_4402 : p19_uge_4402;
      p19_uge_4468 <= p19_data_enable ? p18_uge_4468 : p19_uge_4468;
      p19_uge_4534 <= p19_data_enable ? p18_uge_4534 : p19_uge_4534;
      p19_uge_4600 <= p19_data_enable ? p18_uge_4600 : p19_uge_4600;
      p19_uge_4666 <= p19_data_enable ? p18_uge_4666 : p19_uge_4666;
      p19_uge_4732 <= p19_data_enable ? p18_uge_4732 : p19_uge_4732;
      p19_uge_4798 <= p19_data_enable ? p18_uge_4798 : p19_uge_4798;
      p19_uge_4864 <= p19_data_enable ? p18_uge_4864 : p19_uge_4864;
      p19_uge_4930 <= p19_data_enable ? p18_uge_4930 : p19_uge_4930;
      p19_uge_4996 <= p19_data_enable ? p18_uge_4996 : p19_uge_4996;
      p19_uge_5062 <= p19_data_enable ? p18_uge_5062 : p19_uge_5062;
      p19_uge_5128 <= p19_data_enable ? p18_uge_5128 : p19_uge_5128;
      p19_uge_5194 <= p19_data_enable ? p18_uge_5194 : p19_uge_5194;
      p19_concat_5259 <= p19_data_enable ? concat_5259 : p19_concat_5259;
      p19_uge_5260 <= p19_data_enable ? uge_5260 : p19_uge_5260;
      p19_bit_slice_3986 <= p19_data_enable ? p18_bit_slice_3986 : p19_bit_slice_3986;
      p19_bit_slice_3987 <= p19_data_enable ? p18_bit_slice_3987 : p19_bit_slice_3987;
      p19_bit_slice_3989 <= p19_data_enable ? p18_bit_slice_3989 : p19_bit_slice_3989;
      p19_bit_slice_3990 <= p19_data_enable ? p18_bit_slice_3990 : p19_bit_slice_3990;
      p19_flag_zero <= p19_data_enable ? p18_flag_zero : p19_flag_zero;
      p19_result_sign <= p19_data_enable ? p18_result_sign : p19_result_sign;
      p19_result_exp <= p19_data_enable ? p18_result_exp : p19_result_exp;
      p20_b_fraction <= p20_data_enable ? p19_b_fraction : p20_b_fraction;
      p20_uge_4116 <= p20_data_enable ? p19_uge_4116 : p20_uge_4116;
      p20_b_fractionivisor__1 <= p20_data_enable ? p19_b_fractionivisor__1 : p20_b_fractionivisor__1;
      p20_uge_4124 <= p20_data_enable ? p19_uge_4124 : p20_uge_4124;
      p20_uge_4195 <= p20_data_enable ? p19_uge_4195 : p20_uge_4195;
      p20_uge_4270 <= p20_data_enable ? p19_uge_4270 : p20_uge_4270;
      p20_uge_4336 <= p20_data_enable ? p19_uge_4336 : p20_uge_4336;
      p20_uge_4402 <= p20_data_enable ? p19_uge_4402 : p20_uge_4402;
      p20_uge_4468 <= p20_data_enable ? p19_uge_4468 : p20_uge_4468;
      p20_uge_4534 <= p20_data_enable ? p19_uge_4534 : p20_uge_4534;
      p20_uge_4600 <= p20_data_enable ? p19_uge_4600 : p20_uge_4600;
      p20_uge_4666 <= p20_data_enable ? p19_uge_4666 : p20_uge_4666;
      p20_uge_4732 <= p20_data_enable ? p19_uge_4732 : p20_uge_4732;
      p20_uge_4798 <= p20_data_enable ? p19_uge_4798 : p20_uge_4798;
      p20_uge_4864 <= p20_data_enable ? p19_uge_4864 : p20_uge_4864;
      p20_uge_4930 <= p20_data_enable ? p19_uge_4930 : p20_uge_4930;
      p20_uge_4996 <= p20_data_enable ? p19_uge_4996 : p20_uge_4996;
      p20_uge_5062 <= p20_data_enable ? p19_uge_5062 : p20_uge_5062;
      p20_uge_5128 <= p20_data_enable ? p19_uge_5128 : p20_uge_5128;
      p20_uge_5194 <= p20_data_enable ? p19_uge_5194 : p20_uge_5194;
      p20_uge_5260 <= p20_data_enable ? p19_uge_5260 : p20_uge_5260;
      p20_concat_5325 <= p20_data_enable ? concat_5325 : p20_concat_5325;
      p20_uge_5326 <= p20_data_enable ? uge_5326 : p20_uge_5326;
      p20_bit_slice_3987 <= p20_data_enable ? p19_bit_slice_3987 : p20_bit_slice_3987;
      p20_bit_slice_3989 <= p20_data_enable ? p19_bit_slice_3989 : p20_bit_slice_3989;
      p20_bit_slice_3990 <= p20_data_enable ? p19_bit_slice_3990 : p20_bit_slice_3990;
      p20_flag_zero <= p20_data_enable ? p19_flag_zero : p20_flag_zero;
      p20_result_sign <= p20_data_enable ? p19_result_sign : p20_result_sign;
      p20_result_exp <= p20_data_enable ? p19_result_exp : p20_result_exp;
      p21_b_fraction <= p21_data_enable ? p20_b_fraction : p21_b_fraction;
      p21_uge_4116 <= p21_data_enable ? p20_uge_4116 : p21_uge_4116;
      p21_b_fractionivisor__1 <= p21_data_enable ? p20_b_fractionivisor__1 : p21_b_fractionivisor__1;
      p21_uge_4124 <= p21_data_enable ? p20_uge_4124 : p21_uge_4124;
      p21_uge_4195 <= p21_data_enable ? p20_uge_4195 : p21_uge_4195;
      p21_uge_4270 <= p21_data_enable ? p20_uge_4270 : p21_uge_4270;
      p21_uge_4336 <= p21_data_enable ? p20_uge_4336 : p21_uge_4336;
      p21_uge_4402 <= p21_data_enable ? p20_uge_4402 : p21_uge_4402;
      p21_uge_4468 <= p21_data_enable ? p20_uge_4468 : p21_uge_4468;
      p21_uge_4534 <= p21_data_enable ? p20_uge_4534 : p21_uge_4534;
      p21_uge_4600 <= p21_data_enable ? p20_uge_4600 : p21_uge_4600;
      p21_uge_4666 <= p21_data_enable ? p20_uge_4666 : p21_uge_4666;
      p21_uge_4732 <= p21_data_enable ? p20_uge_4732 : p21_uge_4732;
      p21_uge_4798 <= p21_data_enable ? p20_uge_4798 : p21_uge_4798;
      p21_uge_4864 <= p21_data_enable ? p20_uge_4864 : p21_uge_4864;
      p21_uge_4930 <= p21_data_enable ? p20_uge_4930 : p21_uge_4930;
      p21_uge_4996 <= p21_data_enable ? p20_uge_4996 : p21_uge_4996;
      p21_uge_5062 <= p21_data_enable ? p20_uge_5062 : p21_uge_5062;
      p21_uge_5128 <= p21_data_enable ? p20_uge_5128 : p21_uge_5128;
      p21_uge_5194 <= p21_data_enable ? p20_uge_5194 : p21_uge_5194;
      p21_uge_5260 <= p21_data_enable ? p20_uge_5260 : p21_uge_5260;
      p21_uge_5326 <= p21_data_enable ? p20_uge_5326 : p21_uge_5326;
      p21_concat_5391 <= p21_data_enable ? concat_5391 : p21_concat_5391;
      p21_uge_5392 <= p21_data_enable ? uge_5392 : p21_uge_5392;
      p21_bit_slice_3989 <= p21_data_enable ? p20_bit_slice_3989 : p21_bit_slice_3989;
      p21_bit_slice_3990 <= p21_data_enable ? p20_bit_slice_3990 : p21_bit_slice_3990;
      p21_flag_zero <= p21_data_enable ? p20_flag_zero : p21_flag_zero;
      p21_result_sign <= p21_data_enable ? p20_result_sign : p21_result_sign;
      p21_result_exp <= p21_data_enable ? p20_result_exp : p21_result_exp;
      p22_b_fraction <= p22_data_enable ? p21_b_fraction : p22_b_fraction;
      p22_uge_4116 <= p22_data_enable ? p21_uge_4116 : p22_uge_4116;
      p22_b_fractionivisor__1 <= p22_data_enable ? p21_b_fractionivisor__1 : p22_b_fractionivisor__1;
      p22_uge_4124 <= p22_data_enable ? p21_uge_4124 : p22_uge_4124;
      p22_uge_4195 <= p22_data_enable ? p21_uge_4195 : p22_uge_4195;
      p22_uge_4270 <= p22_data_enable ? p21_uge_4270 : p22_uge_4270;
      p22_uge_4336 <= p22_data_enable ? p21_uge_4336 : p22_uge_4336;
      p22_uge_4402 <= p22_data_enable ? p21_uge_4402 : p22_uge_4402;
      p22_uge_4468 <= p22_data_enable ? p21_uge_4468 : p22_uge_4468;
      p22_uge_4534 <= p22_data_enable ? p21_uge_4534 : p22_uge_4534;
      p22_uge_4600 <= p22_data_enable ? p21_uge_4600 : p22_uge_4600;
      p22_uge_4666 <= p22_data_enable ? p21_uge_4666 : p22_uge_4666;
      p22_uge_4732 <= p22_data_enable ? p21_uge_4732 : p22_uge_4732;
      p22_uge_4798 <= p22_data_enable ? p21_uge_4798 : p22_uge_4798;
      p22_uge_4864 <= p22_data_enable ? p21_uge_4864 : p22_uge_4864;
      p22_uge_4930 <= p22_data_enable ? p21_uge_4930 : p22_uge_4930;
      p22_uge_4996 <= p22_data_enable ? p21_uge_4996 : p22_uge_4996;
      p22_uge_5062 <= p22_data_enable ? p21_uge_5062 : p22_uge_5062;
      p22_uge_5128 <= p22_data_enable ? p21_uge_5128 : p22_uge_5128;
      p22_uge_5194 <= p22_data_enable ? p21_uge_5194 : p22_uge_5194;
      p22_uge_5260 <= p22_data_enable ? p21_uge_5260 : p22_uge_5260;
      p22_uge_5326 <= p22_data_enable ? p21_uge_5326 : p22_uge_5326;
      p22_uge_5392 <= p22_data_enable ? p21_uge_5392 : p22_uge_5392;
      p22_concat_5457 <= p22_data_enable ? concat_5457 : p22_concat_5457;
      p22_uge_5458 <= p22_data_enable ? uge_5458 : p22_uge_5458;
      p22_bit_slice_3990 <= p22_data_enable ? p21_bit_slice_3990 : p22_bit_slice_3990;
      p22_flag_zero <= p22_data_enable ? p21_flag_zero : p22_flag_zero;
      p22_result_sign <= p22_data_enable ? p21_result_sign : p22_result_sign;
      p22_result_exp <= p22_data_enable ? p21_result_exp : p22_result_exp;
      p23_uge_4116 <= p23_data_enable ? p22_uge_4116 : p23_uge_4116;
      p23_uge_4124 <= p23_data_enable ? p22_uge_4124 : p23_uge_4124;
      p23_uge_4195 <= p23_data_enable ? p22_uge_4195 : p23_uge_4195;
      p23_uge_4270 <= p23_data_enable ? p22_uge_4270 : p23_uge_4270;
      p23_uge_4336 <= p23_data_enable ? p22_uge_4336 : p23_uge_4336;
      p23_uge_4402 <= p23_data_enable ? p22_uge_4402 : p23_uge_4402;
      p23_uge_4468 <= p23_data_enable ? p22_uge_4468 : p23_uge_4468;
      p23_uge_4534 <= p23_data_enable ? p22_uge_4534 : p23_uge_4534;
      p23_uge_4600 <= p23_data_enable ? p22_uge_4600 : p23_uge_4600;
      p23_uge_4666 <= p23_data_enable ? p22_uge_4666 : p23_uge_4666;
      p23_uge_4732 <= p23_data_enable ? p22_uge_4732 : p23_uge_4732;
      p23_uge_4798 <= p23_data_enable ? p22_uge_4798 : p23_uge_4798;
      p23_uge_4864 <= p23_data_enable ? p22_uge_4864 : p23_uge_4864;
      p23_uge_4930 <= p23_data_enable ? p22_uge_4930 : p23_uge_4930;
      p23_uge_4996 <= p23_data_enable ? p22_uge_4996 : p23_uge_4996;
      p23_uge_5062 <= p23_data_enable ? p22_uge_5062 : p23_uge_5062;
      p23_uge_5128 <= p23_data_enable ? p22_uge_5128 : p23_uge_5128;
      p23_uge_5194 <= p23_data_enable ? p22_uge_5194 : p23_uge_5194;
      p23_uge_5260 <= p23_data_enable ? p22_uge_5260 : p23_uge_5260;
      p23_uge_5326 <= p23_data_enable ? p22_uge_5326 : p23_uge_5326;
      p23_uge_5392 <= p23_data_enable ? p22_uge_5392 : p23_uge_5392;
      p23_uge_5458 <= p23_data_enable ? p22_uge_5458 : p23_uge_5458;
      p23_flag_zero <= p23_data_enable ? p22_flag_zero : p23_flag_zero;
      p23_q__23_squeezed_portion_0_width_1 <= p23_data_enable ? q__23_squeezed_portion_0_width_1 : p23_q__23_squeezed_portion_0_width_1;
      p23_result_sign <= p23_data_enable ? p22_result_sign : p23_result_sign;
      p23_result_exp <= p23_data_enable ? p22_result_exp : p23_result_exp;
      p0_valid <= p0_enable ? lhs_valid_reg : p0_valid;
      p1_valid <= p1_enable ? p1_stage_done : p1_valid;
      p2_valid <= p2_enable ? p1_valid : p2_valid;
      p3_valid <= p3_enable ? p2_valid : p3_valid;
      p4_valid <= p4_enable ? p3_valid : p4_valid;
      p5_valid <= p5_enable ? p4_valid : p5_valid;
      p6_valid <= p6_enable ? p5_valid : p6_valid;
      p7_valid <= p7_enable ? p6_valid : p7_valid;
      p8_valid <= p8_enable ? p7_valid : p8_valid;
      p9_valid <= p9_enable ? p8_valid : p9_valid;
      p10_valid <= p10_enable ? p9_valid : p10_valid;
      p11_valid <= p11_enable ? p10_valid : p11_valid;
      p12_valid <= p12_enable ? p11_valid : p12_valid;
      p13_valid <= p13_enable ? p12_valid : p13_valid;
      p14_valid <= p14_enable ? p13_valid : p14_valid;
      p15_valid <= p15_enable ? p14_valid : p15_valid;
      p16_valid <= p16_enable ? p15_valid : p16_valid;
      p17_valid <= p17_enable ? p16_valid : p17_valid;
      p18_valid <= p18_enable ? p17_valid : p18_valid;
      p19_valid <= p19_enable ? p18_valid : p19_valid;
      p20_valid <= p20_enable ? p19_valid : p20_valid;
      p21_valid <= p21_enable ? p20_valid : p21_valid;
      p22_valid <= p22_enable ? p21_valid : p22_valid;
      p23_valid <= p23_enable ? p22_valid : p23_valid;
      p24_valid <= p24_enable ? p24_stage_done : p24_valid;
      p25_valid <= p25_enable ? p24_valid : p25_valid;
      p26_valid <= p26_enable ? p25_valid : p26_valid;
      p27_valid <= p27_enable ? p26_valid : p27_valid;
      p28_valid <= p28_enable ? p27_valid : p28_valid;
      p29_valid <= p29_enable ? p28_valid : p29_valid;
      p30_valid <= p30_enable ? p29_valid : p30_valid;
      lhs_reg <= lhs_load_en ? lhs : lhs_reg;
      lhs_valid_reg <= lhs_valid_load_en ? lhs_valid : lhs_valid_reg;
      rhs_reg <= rhs_load_en ? rhs : rhs_reg;
      rhs_valid_reg <= rhs_valid_load_en ? rhs_valid : rhs_valid_reg;
      result_reg <= result_load_en ? sum : result_reg;
      result_valid_reg <= result_valid_load_en ? p23_valid : result_valid_reg;
    end
  end
  assign result = result_reg;
  assign result_valid = result_valid_reg;
  assign lhs_ready = lhs_load_en;
  assign rhs_ready = rhs_load_en;
endmodule
module xls_divsi32(
  input wire clk,
  input wire rst,
  input wire [31:0] lhs,
  input wire lhs_valid,
  input wire [31:0] rhs,
  input wire rhs_valid,
  input wire result_ready,
  output wire [31:0] result,
  output wire result_valid,
  output wire lhs_ready,
  output wire rhs_ready
);
  reg p0_sign_a;
  reg [31:0] p0_b;
  reg p0_bit_slice_6525;
  reg p0_bit_slice_6526;
  reg p0_bit_slice_6527;
  reg p0_bit_slice_6528;
  reg p0_bit_slice_6529;
  reg p0_bit_slice_6530;
  reg p0_bit_slice_6531;
  reg p0_bit_slice_6532;
  reg p0_bit_slice_6533;
  reg p0_bit_slice_6534;
  reg p0_bit_slice_6535;
  reg p0_bit_slice_6536;
  reg p0_bit_slice_6537;
  reg p0_bit_slice_6538;
  reg p0_bit_slice_6539;
  reg p0_bit_slice_6540;
  reg p0_bit_slice_6541;
  reg p0_bit_slice_6542;
  reg p0_bit_slice_6543;
  reg p0_bit_slice_6544;
  reg p0_bit_slice_6545;
  reg p0_bit_slice_6546;
  reg p0_bit_slice_6547;
  reg p0_bit_slice_6548;
  reg p0_bit_slice_6549;
  reg p0_bit_slice_6550;
  reg p0_bit_slice_6551;
  reg p0_bit_slice_6552;
  reg p0_bit_slice_6553;
  reg p0_bit_slice_6554;
  reg p0_bit_slice_6555;
  reg [31:0] p1_b;
  reg p1_uge_6629;
  reg [32:0] p1_bivisor__1;
  reg [31:0] p1_concat_6636;
  reg p1_uge_6637;
  reg p1_bit_slice_6526;
  reg p1_bit_slice_6527;
  reg p1_bit_slice_6528;
  reg p1_bit_slice_6529;
  reg p1_bit_slice_6530;
  reg p1_bit_slice_6531;
  reg p1_bit_slice_6532;
  reg p1_bit_slice_6533;
  reg p1_bit_slice_6534;
  reg p1_bit_slice_6535;
  reg p1_bit_slice_6536;
  reg p1_bit_slice_6537;
  reg p1_bit_slice_6538;
  reg p1_bit_slice_6539;
  reg p1_bit_slice_6540;
  reg p1_bit_slice_6541;
  reg p1_bit_slice_6542;
  reg p1_bit_slice_6543;
  reg p1_bit_slice_6544;
  reg p1_bit_slice_6545;
  reg p1_bit_slice_6546;
  reg p1_bit_slice_6547;
  reg p1_bit_slice_6548;
  reg p1_bit_slice_6549;
  reg p1_bit_slice_6550;
  reg p1_bit_slice_6551;
  reg p1_bit_slice_6552;
  reg p1_bit_slice_6553;
  reg p1_bit_slice_6554;
  reg p1_bit_slice_6555;
  reg p1_negated;
  reg [31:0] p2_b;
  reg p2_uge_6629;
  reg [32:0] p2_bivisor__1;
  reg p2_uge_6637;
  reg [31:0] p2_concat_6718;
  reg p2_uge_6719;
  reg [31:0] p2_sub_6720;
  reg p2_bit_slice_6527;
  reg p2_bit_slice_6528;
  reg p2_bit_slice_6529;
  reg p2_bit_slice_6530;
  reg p2_bit_slice_6531;
  reg p2_bit_slice_6532;
  reg p2_bit_slice_6533;
  reg p2_bit_slice_6534;
  reg p2_bit_slice_6535;
  reg p2_bit_slice_6536;
  reg p2_bit_slice_6537;
  reg p2_bit_slice_6538;
  reg p2_bit_slice_6539;
  reg p2_bit_slice_6540;
  reg p2_bit_slice_6541;
  reg p2_bit_slice_6542;
  reg p2_bit_slice_6543;
  reg p2_bit_slice_6544;
  reg p2_bit_slice_6545;
  reg p2_bit_slice_6546;
  reg p2_bit_slice_6547;
  reg p2_bit_slice_6548;
  reg p2_bit_slice_6549;
  reg p2_bit_slice_6550;
  reg p2_bit_slice_6551;
  reg p2_bit_slice_6552;
  reg p2_bit_slice_6553;
  reg p2_bit_slice_6554;
  reg p2_bit_slice_6555;
  reg p2_negated;
  reg [31:0] p3_b;
  reg p3_uge_6629;
  reg [32:0] p3_bivisor__1;
  reg p3_uge_6637;
  reg p3_uge_6719;
  reg p3_uge_6801;
  reg [31:0] p3_r__68;
  reg p3_bit_slice_6528;
  reg p3_bit_slice_6529;
  reg p3_bit_slice_6530;
  reg p3_bit_slice_6531;
  reg p3_bit_slice_6532;
  reg p3_bit_slice_6533;
  reg p3_bit_slice_6534;
  reg p3_bit_slice_6535;
  reg p3_bit_slice_6536;
  reg p3_bit_slice_6537;
  reg p3_bit_slice_6538;
  reg p3_bit_slice_6539;
  reg p3_bit_slice_6540;
  reg p3_bit_slice_6541;
  reg p3_bit_slice_6542;
  reg p3_bit_slice_6543;
  reg p3_bit_slice_6544;
  reg p3_bit_slice_6545;
  reg p3_bit_slice_6546;
  reg p3_bit_slice_6547;
  reg p3_bit_slice_6548;
  reg p3_bit_slice_6549;
  reg p3_bit_slice_6550;
  reg p3_bit_slice_6551;
  reg p3_bit_slice_6552;
  reg p3_bit_slice_6553;
  reg p3_bit_slice_6554;
  reg p3_bit_slice_6555;
  reg p3_negated;
  reg [31:0] p4_b;
  reg p4_uge_6629;
  reg [32:0] p4_bivisor__1;
  reg p4_uge_6637;
  reg p4_uge_6719;
  reg p4_uge_6801;
  reg p4_uge_6881;
  reg [31:0] p4_r__69;
  reg p4_bit_slice_6529;
  reg [30:0] p4_bit_slice_6884;
  reg p4_bit_slice_6530;
  reg p4_bit_slice_6531;
  reg p4_bit_slice_6532;
  reg p4_bit_slice_6533;
  reg p4_bit_slice_6534;
  reg p4_bit_slice_6535;
  reg p4_bit_slice_6536;
  reg p4_bit_slice_6537;
  reg p4_bit_slice_6538;
  reg p4_bit_slice_6539;
  reg p4_bit_slice_6540;
  reg p4_bit_slice_6541;
  reg p4_bit_slice_6542;
  reg p4_bit_slice_6543;
  reg p4_bit_slice_6544;
  reg p4_bit_slice_6545;
  reg p4_bit_slice_6546;
  reg p4_bit_slice_6547;
  reg p4_bit_slice_6548;
  reg p4_bit_slice_6549;
  reg p4_bit_slice_6550;
  reg p4_bit_slice_6551;
  reg p4_bit_slice_6552;
  reg p4_bit_slice_6553;
  reg p4_bit_slice_6554;
  reg p4_bit_slice_6555;
  reg p4_negated;
  reg [31:0] p5_b;
  reg p5_uge_6629;
  reg [32:0] p5_bivisor__1;
  reg p5_uge_6637;
  reg p5_uge_6719;
  reg p5_uge_6801;
  reg p5_uge_6881;
  reg p5_uge_6963;
  reg [31:0] p5_concat_6968;
  reg p5_uge_6969;
  reg p5_bit_slice_6531;
  reg p5_bit_slice_6532;
  reg p5_bit_slice_6533;
  reg p5_bit_slice_6534;
  reg p5_bit_slice_6535;
  reg p5_bit_slice_6536;
  reg p5_bit_slice_6537;
  reg p5_bit_slice_6538;
  reg p5_bit_slice_6539;
  reg p5_bit_slice_6540;
  reg p5_bit_slice_6541;
  reg p5_bit_slice_6542;
  reg p5_bit_slice_6543;
  reg p5_bit_slice_6544;
  reg p5_bit_slice_6545;
  reg p5_bit_slice_6546;
  reg p5_bit_slice_6547;
  reg p5_bit_slice_6548;
  reg p5_bit_slice_6549;
  reg p5_bit_slice_6550;
  reg p5_bit_slice_6551;
  reg p5_bit_slice_6552;
  reg p5_bit_slice_6553;
  reg p5_bit_slice_6554;
  reg p5_bit_slice_6555;
  reg p5_negated;
  reg [31:0] p6_b;
  reg p6_uge_6629;
  reg [32:0] p6_bivisor__1;
  reg p6_uge_6637;
  reg p6_uge_6719;
  reg p6_uge_6801;
  reg p6_uge_6881;
  reg p6_uge_6963;
  reg p6_uge_6969;
  reg [31:0] p6_concat_7048;
  reg p6_uge_7049;
  reg [31:0] p6_sub_7050;
  reg p6_bit_slice_6532;
  reg p6_bit_slice_6533;
  reg p6_bit_slice_6534;
  reg p6_bit_slice_6535;
  reg p6_bit_slice_6536;
  reg p6_bit_slice_6537;
  reg p6_bit_slice_6538;
  reg p6_bit_slice_6539;
  reg p6_bit_slice_6540;
  reg p6_bit_slice_6541;
  reg p6_bit_slice_6542;
  reg p6_bit_slice_6543;
  reg p6_bit_slice_6544;
  reg p6_bit_slice_6545;
  reg p6_bit_slice_6546;
  reg p6_bit_slice_6547;
  reg p6_bit_slice_6548;
  reg p6_bit_slice_6549;
  reg p6_bit_slice_6550;
  reg p6_bit_slice_6551;
  reg p6_bit_slice_6552;
  reg p6_bit_slice_6553;
  reg p6_bit_slice_6554;
  reg p6_bit_slice_6555;
  reg p6_negated;
  reg [31:0] p7_b;
  reg p7_uge_6629;
  reg [32:0] p7_bivisor__1;
  reg p7_uge_6637;
  reg p7_uge_6719;
  reg p7_uge_6801;
  reg p7_uge_6881;
  reg p7_uge_6963;
  reg p7_uge_6969;
  reg p7_uge_7049;
  reg p7_uge_7131;
  reg [31:0] p7_r__73;
  reg p7_bit_slice_6533;
  reg p7_bit_slice_6534;
  reg p7_bit_slice_6535;
  reg p7_bit_slice_6536;
  reg p7_bit_slice_6537;
  reg p7_bit_slice_6538;
  reg p7_bit_slice_6539;
  reg p7_bit_slice_6540;
  reg p7_bit_slice_6541;
  reg p7_bit_slice_6542;
  reg p7_bit_slice_6543;
  reg p7_bit_slice_6544;
  reg p7_bit_slice_6545;
  reg p7_bit_slice_6546;
  reg p7_bit_slice_6547;
  reg p7_bit_slice_6548;
  reg p7_bit_slice_6549;
  reg p7_bit_slice_6550;
  reg p7_bit_slice_6551;
  reg p7_bit_slice_6552;
  reg p7_bit_slice_6553;
  reg p7_bit_slice_6554;
  reg p7_bit_slice_6555;
  reg p7_negated;
  reg [31:0] p8_b;
  reg p8_uge_6629;
  reg [32:0] p8_bivisor__1;
  reg p8_uge_6637;
  reg p8_uge_6719;
  reg p8_uge_6801;
  reg p8_uge_6881;
  reg p8_uge_6963;
  reg p8_uge_6969;
  reg p8_uge_7049;
  reg p8_uge_7131;
  reg p8_uge_7211;
  reg [31:0] p8_r__74;
  reg p8_bit_slice_6534;
  reg [30:0] p8_bit_slice_7214;
  reg p8_bit_slice_6535;
  reg p8_bit_slice_6536;
  reg p8_bit_slice_6537;
  reg p8_bit_slice_6538;
  reg p8_bit_slice_6539;
  reg p8_bit_slice_6540;
  reg p8_bit_slice_6541;
  reg p8_bit_slice_6542;
  reg p8_bit_slice_6543;
  reg p8_bit_slice_6544;
  reg p8_bit_slice_6545;
  reg p8_bit_slice_6546;
  reg p8_bit_slice_6547;
  reg p8_bit_slice_6548;
  reg p8_bit_slice_6549;
  reg p8_bit_slice_6550;
  reg p8_bit_slice_6551;
  reg p8_bit_slice_6552;
  reg p8_bit_slice_6553;
  reg p8_bit_slice_6554;
  reg p8_bit_slice_6555;
  reg p8_negated;
  reg [31:0] p9_b;
  reg p9_uge_6629;
  reg [32:0] p9_bivisor__1;
  reg p9_uge_6637;
  reg p9_uge_6719;
  reg p9_uge_6801;
  reg p9_uge_6881;
  reg p9_uge_6963;
  reg p9_uge_6969;
  reg p9_uge_7049;
  reg p9_uge_7131;
  reg p9_uge_7211;
  reg p9_uge_7293;
  reg [31:0] p9_concat_7298;
  reg p9_uge_7299;
  reg p9_bit_slice_6536;
  reg p9_bit_slice_6537;
  reg p9_bit_slice_6538;
  reg p9_bit_slice_6539;
  reg p9_bit_slice_6540;
  reg p9_bit_slice_6541;
  reg p9_bit_slice_6542;
  reg p9_bit_slice_6543;
  reg p9_bit_slice_6544;
  reg p9_bit_slice_6545;
  reg p9_bit_slice_6546;
  reg p9_bit_slice_6547;
  reg p9_bit_slice_6548;
  reg p9_bit_slice_6549;
  reg p9_bit_slice_6550;
  reg p9_bit_slice_6551;
  reg p9_bit_slice_6552;
  reg p9_bit_slice_6553;
  reg p9_bit_slice_6554;
  reg p9_bit_slice_6555;
  reg p9_negated;
  reg [31:0] p10_b;
  reg p10_uge_6629;
  reg [32:0] p10_bivisor__1;
  reg p10_uge_6637;
  reg p10_uge_6719;
  reg p10_uge_6801;
  reg p10_uge_6881;
  reg p10_uge_6963;
  reg p10_uge_6969;
  reg p10_uge_7049;
  reg p10_uge_7131;
  reg p10_uge_7211;
  reg p10_uge_7293;
  reg p10_uge_7299;
  reg [31:0] p10_concat_7378;
  reg p10_uge_7379;
  reg [31:0] p10_sub_7380;
  reg p10_bit_slice_6537;
  reg p10_bit_slice_6538;
  reg p10_bit_slice_6539;
  reg p10_bit_slice_6540;
  reg p10_bit_slice_6541;
  reg p10_bit_slice_6542;
  reg p10_bit_slice_6543;
  reg p10_bit_slice_6544;
  reg p10_bit_slice_6545;
  reg p10_bit_slice_6546;
  reg p10_bit_slice_6547;
  reg p10_bit_slice_6548;
  reg p10_bit_slice_6549;
  reg p10_bit_slice_6550;
  reg p10_bit_slice_6551;
  reg p10_bit_slice_6552;
  reg p10_bit_slice_6553;
  reg p10_bit_slice_6554;
  reg p10_bit_slice_6555;
  reg p10_negated;
  reg [31:0] p11_b;
  reg p11_uge_6629;
  reg [32:0] p11_bivisor__1;
  reg p11_uge_6637;
  reg p11_uge_6719;
  reg p11_uge_6801;
  reg p11_uge_6881;
  reg p11_uge_6963;
  reg p11_uge_6969;
  reg p11_uge_7049;
  reg p11_uge_7131;
  reg p11_uge_7211;
  reg p11_uge_7293;
  reg p11_uge_7299;
  reg p11_uge_7379;
  reg p11_uge_7461;
  reg [31:0] p11_r__78;
  reg p11_bit_slice_6538;
  reg p11_bit_slice_6539;
  reg p11_bit_slice_6540;
  reg p11_bit_slice_6541;
  reg p11_bit_slice_6542;
  reg p11_bit_slice_6543;
  reg p11_bit_slice_6544;
  reg p11_bit_slice_6545;
  reg p11_bit_slice_6546;
  reg p11_bit_slice_6547;
  reg p11_bit_slice_6548;
  reg p11_bit_slice_6549;
  reg p11_bit_slice_6550;
  reg p11_bit_slice_6551;
  reg p11_bit_slice_6552;
  reg p11_bit_slice_6553;
  reg p11_bit_slice_6554;
  reg p11_bit_slice_6555;
  reg p11_negated;
  reg [31:0] p12_b;
  reg p12_uge_6629;
  reg [32:0] p12_bivisor__1;
  reg p12_uge_6637;
  reg p12_uge_6719;
  reg p12_uge_6801;
  reg p12_uge_6881;
  reg p12_uge_6963;
  reg p12_uge_6969;
  reg p12_uge_7049;
  reg p12_uge_7131;
  reg p12_uge_7211;
  reg p12_uge_7293;
  reg p12_uge_7299;
  reg p12_uge_7379;
  reg p12_uge_7461;
  reg p12_uge_7541;
  reg [31:0] p12_r__79;
  reg p12_bit_slice_6539;
  reg [30:0] p12_bit_slice_7544;
  reg p12_bit_slice_6540;
  reg p12_bit_slice_6541;
  reg p12_bit_slice_6542;
  reg p12_bit_slice_6543;
  reg p12_bit_slice_6544;
  reg p12_bit_slice_6545;
  reg p12_bit_slice_6546;
  reg p12_bit_slice_6547;
  reg p12_bit_slice_6548;
  reg p12_bit_slice_6549;
  reg p12_bit_slice_6550;
  reg p12_bit_slice_6551;
  reg p12_bit_slice_6552;
  reg p12_bit_slice_6553;
  reg p12_bit_slice_6554;
  reg p12_bit_slice_6555;
  reg p12_negated;
  reg [31:0] p13_b;
  reg p13_uge_6629;
  reg [32:0] p13_bivisor__1;
  reg p13_uge_6637;
  reg p13_uge_6719;
  reg p13_uge_6801;
  reg p13_uge_6881;
  reg p13_uge_6963;
  reg p13_uge_6969;
  reg p13_uge_7049;
  reg p13_uge_7131;
  reg p13_uge_7211;
  reg p13_uge_7293;
  reg p13_uge_7299;
  reg p13_uge_7379;
  reg p13_uge_7461;
  reg p13_uge_7541;
  reg p13_uge_7623;
  reg [31:0] p13_concat_7628;
  reg p13_uge_7629;
  reg p13_bit_slice_6541;
  reg p13_bit_slice_6542;
  reg p13_bit_slice_6543;
  reg p13_bit_slice_6544;
  reg p13_bit_slice_6545;
  reg p13_bit_slice_6546;
  reg p13_bit_slice_6547;
  reg p13_bit_slice_6548;
  reg p13_bit_slice_6549;
  reg p13_bit_slice_6550;
  reg p13_bit_slice_6551;
  reg p13_bit_slice_6552;
  reg p13_bit_slice_6553;
  reg p13_bit_slice_6554;
  reg p13_bit_slice_6555;
  reg p13_negated;
  reg [31:0] p14_b;
  reg p14_uge_6629;
  reg [32:0] p14_bivisor__1;
  reg p14_uge_6637;
  reg p14_uge_6719;
  reg p14_uge_6801;
  reg p14_uge_6881;
  reg p14_uge_6963;
  reg p14_uge_6969;
  reg p14_uge_7049;
  reg p14_uge_7131;
  reg p14_uge_7211;
  reg p14_uge_7293;
  reg p14_uge_7299;
  reg p14_uge_7379;
  reg p14_uge_7461;
  reg p14_uge_7541;
  reg p14_uge_7623;
  reg p14_uge_7629;
  reg [31:0] p14_concat_7708;
  reg p14_uge_7709;
  reg [31:0] p14_sub_7710;
  reg p14_bit_slice_6542;
  reg p14_bit_slice_6543;
  reg p14_bit_slice_6544;
  reg p14_bit_slice_6545;
  reg p14_bit_slice_6546;
  reg p14_bit_slice_6547;
  reg p14_bit_slice_6548;
  reg p14_bit_slice_6549;
  reg p14_bit_slice_6550;
  reg p14_bit_slice_6551;
  reg p14_bit_slice_6552;
  reg p14_bit_slice_6553;
  reg p14_bit_slice_6554;
  reg p14_bit_slice_6555;
  reg p14_negated;
  reg [31:0] p15_b;
  reg p15_uge_6629;
  reg [32:0] p15_bivisor__1;
  reg p15_uge_6637;
  reg p15_uge_6719;
  reg p15_uge_6801;
  reg p15_uge_6881;
  reg p15_uge_6963;
  reg p15_uge_6969;
  reg p15_uge_7049;
  reg p15_uge_7131;
  reg p15_uge_7211;
  reg p15_uge_7293;
  reg p15_uge_7299;
  reg p15_uge_7379;
  reg p15_uge_7461;
  reg p15_uge_7541;
  reg p15_uge_7623;
  reg p15_uge_7629;
  reg p15_uge_7709;
  reg p15_uge_7791;
  reg [31:0] p15_r__83;
  reg p15_bit_slice_6543;
  reg p15_bit_slice_6544;
  reg p15_bit_slice_6545;
  reg p15_bit_slice_6546;
  reg p15_bit_slice_6547;
  reg p15_bit_slice_6548;
  reg p15_bit_slice_6549;
  reg p15_bit_slice_6550;
  reg p15_bit_slice_6551;
  reg p15_bit_slice_6552;
  reg p15_bit_slice_6553;
  reg p15_bit_slice_6554;
  reg p15_bit_slice_6555;
  reg p15_negated;
  reg [31:0] p16_b;
  reg p16_uge_6629;
  reg [32:0] p16_bivisor__1;
  reg p16_uge_6637;
  reg p16_uge_6719;
  reg p16_uge_6801;
  reg p16_uge_6881;
  reg p16_uge_6963;
  reg p16_uge_6969;
  reg p16_uge_7049;
  reg p16_uge_7131;
  reg p16_uge_7211;
  reg p16_uge_7293;
  reg p16_uge_7299;
  reg p16_uge_7379;
  reg p16_uge_7461;
  reg p16_uge_7541;
  reg p16_uge_7623;
  reg p16_uge_7629;
  reg p16_uge_7709;
  reg p16_uge_7791;
  reg p16_uge_7871;
  reg [31:0] p16_r__84;
  reg p16_bit_slice_6544;
  reg [30:0] p16_bit_slice_7874;
  reg p16_bit_slice_6545;
  reg p16_bit_slice_6546;
  reg p16_bit_slice_6547;
  reg p16_bit_slice_6548;
  reg p16_bit_slice_6549;
  reg p16_bit_slice_6550;
  reg p16_bit_slice_6551;
  reg p16_bit_slice_6552;
  reg p16_bit_slice_6553;
  reg p16_bit_slice_6554;
  reg p16_bit_slice_6555;
  reg p16_negated;
  reg [31:0] p17_b;
  reg p17_uge_6629;
  reg [32:0] p17_bivisor__1;
  reg p17_uge_6637;
  reg p17_uge_6719;
  reg p17_uge_6801;
  reg p17_uge_6881;
  reg p17_uge_6963;
  reg p17_uge_6969;
  reg p17_uge_7049;
  reg p17_uge_7131;
  reg p17_uge_7211;
  reg p17_uge_7293;
  reg p17_uge_7299;
  reg p17_uge_7379;
  reg p17_uge_7461;
  reg p17_uge_7541;
  reg p17_uge_7623;
  reg p17_uge_7629;
  reg p17_uge_7709;
  reg p17_uge_7791;
  reg p17_uge_7871;
  reg p17_uge_7953;
  reg [31:0] p17_concat_7958;
  reg p17_uge_7959;
  reg p17_bit_slice_6546;
  reg p17_bit_slice_6547;
  reg p17_bit_slice_6548;
  reg p17_bit_slice_6549;
  reg p17_bit_slice_6550;
  reg p17_bit_slice_6551;
  reg p17_bit_slice_6552;
  reg p17_bit_slice_6553;
  reg p17_bit_slice_6554;
  reg p17_bit_slice_6555;
  reg p17_negated;
  reg [31:0] p18_b;
  reg p18_uge_6629;
  reg [32:0] p18_bivisor__1;
  reg p18_uge_6637;
  reg p18_uge_6719;
  reg p18_uge_6801;
  reg p18_uge_6881;
  reg p18_uge_6963;
  reg p18_uge_6969;
  reg p18_uge_7049;
  reg p18_uge_7131;
  reg p18_uge_7211;
  reg p18_uge_7293;
  reg p18_uge_7299;
  reg p18_uge_7379;
  reg p18_uge_7461;
  reg p18_uge_7541;
  reg p18_uge_7623;
  reg p18_uge_7629;
  reg p18_uge_7709;
  reg p18_uge_7791;
  reg p18_uge_7871;
  reg p18_uge_7953;
  reg p18_uge_7959;
  reg [31:0] p18_concat_8038;
  reg p18_uge_8039;
  reg [31:0] p18_sub_8040;
  reg p18_bit_slice_6547;
  reg p18_bit_slice_6548;
  reg p18_bit_slice_6549;
  reg p18_bit_slice_6550;
  reg p18_bit_slice_6551;
  reg p18_bit_slice_6552;
  reg p18_bit_slice_6553;
  reg p18_bit_slice_6554;
  reg p18_bit_slice_6555;
  reg p18_negated;
  reg [31:0] p19_b;
  reg p19_uge_6629;
  reg [32:0] p19_bivisor__1;
  reg p19_uge_6637;
  reg p19_uge_6719;
  reg p19_uge_6801;
  reg p19_uge_6881;
  reg p19_uge_6963;
  reg p19_uge_6969;
  reg p19_uge_7049;
  reg p19_uge_7131;
  reg p19_uge_7211;
  reg p19_uge_7293;
  reg p19_uge_7299;
  reg p19_uge_7379;
  reg p19_uge_7461;
  reg p19_uge_7541;
  reg p19_uge_7623;
  reg p19_uge_7629;
  reg p19_uge_7709;
  reg p19_uge_7791;
  reg p19_uge_7871;
  reg p19_uge_7953;
  reg p19_uge_7959;
  reg p19_uge_8039;
  reg p19_uge_8121;
  reg [31:0] p19_r__88;
  reg p19_bit_slice_6548;
  reg p19_bit_slice_6549;
  reg p19_bit_slice_6550;
  reg p19_bit_slice_6551;
  reg p19_bit_slice_6552;
  reg p19_bit_slice_6553;
  reg p19_bit_slice_6554;
  reg p19_bit_slice_6555;
  reg p19_negated;
  reg [31:0] p20_b;
  reg p20_uge_6629;
  reg [32:0] p20_bivisor__1;
  reg p20_uge_6637;
  reg p20_uge_6719;
  reg p20_uge_6801;
  reg p20_uge_6881;
  reg p20_uge_6963;
  reg p20_uge_6969;
  reg p20_uge_7049;
  reg p20_uge_7131;
  reg p20_uge_7211;
  reg p20_uge_7293;
  reg p20_uge_7299;
  reg p20_uge_7379;
  reg p20_uge_7461;
  reg p20_uge_7541;
  reg p20_uge_7623;
  reg p20_uge_7629;
  reg p20_uge_7709;
  reg p20_uge_7791;
  reg p20_uge_7871;
  reg p20_uge_7953;
  reg p20_uge_7959;
  reg p20_uge_8039;
  reg p20_uge_8121;
  reg p20_uge_8201;
  reg [31:0] p20_r__89;
  reg p20_bit_slice_6549;
  reg [30:0] p20_bit_slice_8204;
  reg p20_bit_slice_6550;
  reg p20_bit_slice_6551;
  reg p20_bit_slice_6552;
  reg p20_bit_slice_6553;
  reg p20_bit_slice_6554;
  reg p20_bit_slice_6555;
  reg p20_negated;
  reg [31:0] p21_b;
  reg p21_uge_6629;
  reg [32:0] p21_bivisor__1;
  reg p21_uge_6637;
  reg p21_uge_6719;
  reg p21_uge_6801;
  reg p21_uge_6881;
  reg p21_uge_6963;
  reg p21_uge_6969;
  reg p21_uge_7049;
  reg p21_uge_7131;
  reg p21_uge_7211;
  reg p21_uge_7293;
  reg p21_uge_7299;
  reg p21_uge_7379;
  reg p21_uge_7461;
  reg p21_uge_7541;
  reg p21_uge_7623;
  reg p21_uge_7629;
  reg p21_uge_7709;
  reg p21_uge_7791;
  reg p21_uge_7871;
  reg p21_uge_7953;
  reg p21_uge_7959;
  reg p21_uge_8039;
  reg p21_uge_8121;
  reg p21_uge_8201;
  reg p21_uge_8283;
  reg [31:0] p21_concat_8288;
  reg p21_uge_8289;
  reg p21_bit_slice_6551;
  reg p21_bit_slice_6552;
  reg p21_bit_slice_6553;
  reg p21_bit_slice_6554;
  reg p21_bit_slice_6555;
  reg p21_negated;
  reg [31:0] p22_b;
  reg p22_uge_6629;
  reg [32:0] p22_bivisor__1;
  reg p22_uge_6637;
  reg p22_uge_6719;
  reg p22_uge_6801;
  reg p22_uge_6881;
  reg p22_uge_6963;
  reg p22_uge_6969;
  reg p22_uge_7049;
  reg p22_uge_7131;
  reg p22_uge_7211;
  reg p22_uge_7293;
  reg p22_uge_7299;
  reg p22_uge_7379;
  reg p22_uge_7461;
  reg p22_uge_7541;
  reg p22_uge_7623;
  reg p22_uge_7629;
  reg p22_uge_7709;
  reg p22_uge_7791;
  reg p22_uge_7871;
  reg p22_uge_7953;
  reg p22_uge_7959;
  reg p22_uge_8039;
  reg p22_uge_8121;
  reg p22_uge_8201;
  reg p22_uge_8283;
  reg p22_uge_8289;
  reg [31:0] p22_concat_8368;
  reg p22_uge_8369;
  reg [31:0] p22_sub_8370;
  reg p22_bit_slice_6552;
  reg p22_bit_slice_6553;
  reg p22_bit_slice_6554;
  reg p22_bit_slice_6555;
  reg p22_negated;
  reg [31:0] p23_b;
  reg p23_uge_6629;
  reg [32:0] p23_bivisor__1;
  reg p23_uge_6637;
  reg p23_uge_6719;
  reg p23_uge_6801;
  reg p23_uge_6881;
  reg p23_uge_6963;
  reg p23_uge_6969;
  reg p23_uge_7049;
  reg p23_uge_7131;
  reg p23_uge_7211;
  reg p23_uge_7293;
  reg p23_uge_7299;
  reg p23_uge_7379;
  reg p23_uge_7461;
  reg p23_uge_7541;
  reg p23_uge_7623;
  reg p23_uge_7629;
  reg p23_uge_7709;
  reg p23_uge_7791;
  reg p23_uge_7871;
  reg p23_uge_7953;
  reg p23_uge_7959;
  reg p23_uge_8039;
  reg p23_uge_8121;
  reg p23_uge_8201;
  reg p23_uge_8283;
  reg p23_uge_8289;
  reg p23_uge_8369;
  reg p23_uge_8451;
  reg [31:0] p23_r__93;
  reg p23_bit_slice_6553;
  reg p23_bit_slice_6554;
  reg p23_bit_slice_6555;
  reg p23_negated;
  reg [31:0] p24_b;
  reg p24_uge_6629;
  reg [32:0] p24_bivisor__1;
  reg p24_uge_6637;
  reg p24_uge_6719;
  reg p24_uge_6801;
  reg p24_uge_6881;
  reg p24_uge_6963;
  reg p24_uge_6969;
  reg p24_uge_7049;
  reg p24_uge_7131;
  reg p24_uge_7211;
  reg p24_uge_7293;
  reg p24_uge_7299;
  reg p24_uge_7379;
  reg p24_uge_7461;
  reg p24_uge_7541;
  reg p24_uge_7623;
  reg p24_uge_7629;
  reg p24_uge_7709;
  reg p24_uge_7791;
  reg p24_uge_7871;
  reg p24_uge_7953;
  reg p24_uge_7959;
  reg p24_uge_8039;
  reg p24_uge_8121;
  reg p24_uge_8201;
  reg p24_uge_8283;
  reg p24_uge_8289;
  reg p24_uge_8369;
  reg p24_uge_8451;
  reg p24_uge_8531;
  reg [31:0] p24_r__94;
  reg p24_bit_slice_6554;
  reg [30:0] p24_bit_slice_8534;
  reg p24_bit_slice_6555;
  reg p24_negated;
  reg p25_uge_6629;
  reg p25_uge_6637;
  reg p25_uge_6719;
  reg p25_uge_6801;
  reg p25_uge_6881;
  reg p25_uge_6963;
  reg p25_uge_6969;
  reg p25_uge_7049;
  reg p25_uge_7131;
  reg p25_uge_7211;
  reg p25_uge_7293;
  reg p25_uge_7299;
  reg p25_uge_7379;
  reg p25_uge_7461;
  reg p25_uge_7541;
  reg p25_uge_7623;
  reg p25_uge_7629;
  reg p25_uge_7709;
  reg p25_uge_7791;
  reg p25_uge_7871;
  reg p25_uge_7953;
  reg p25_uge_7959;
  reg p25_uge_8039;
  reg p25_uge_8121;
  reg p25_uge_8201;
  reg p25_uge_8283;
  reg p25_uge_8289;
  reg p25_uge_8369;
  reg p25_uge_8451;
  reg p25_uge_8531;
  reg p25_uge_8613;
  reg p25_q__32_squeezed_portion_0_width_1;
  reg p25_negated;
  reg p0_valid;
  reg p1_valid;
  reg p2_valid;
  reg p3_valid;
  reg p4_valid;
  reg p5_valid;
  reg p6_valid;
  reg p7_valid;
  reg p8_valid;
  reg p9_valid;
  reg p10_valid;
  reg p11_valid;
  reg p12_valid;
  reg p13_valid;
  reg p14_valid;
  reg p15_valid;
  reg p16_valid;
  reg p17_valid;
  reg p18_valid;
  reg p19_valid;
  reg p20_valid;
  reg p21_valid;
  reg p22_valid;
  reg p23_valid;
  reg p24_valid;
  reg p25_valid;
  reg p26_valid;
  reg p27_valid;
  reg p28_valid;
  reg p29_valid;
  reg p30_valid;
  reg [31:0] lhs_reg;
  reg lhs_valid_reg;
  reg [31:0] rhs_reg;
  reg rhs_valid_reg;
  reg [31:0] result_reg;
  reg result_valid_reg;
  wire result_valid_inv;
  wire result_valid_load_en;
  wire result_load_en;
  wire p26_stage_done;
  wire p26_not_valid;
  wire p25_enable;
  wire p25_data_enable;
  wire p25_not_valid;
  wire p24_enable;
  wire p24_data_enable;
  wire p24_not_valid;
  wire p23_enable;
  wire p23_data_enable;
  wire p23_not_valid;
  wire p22_enable;
  wire p22_data_enable;
  wire p22_not_valid;
  wire p21_enable;
  wire p21_data_enable;
  wire p21_not_valid;
  wire p20_enable;
  wire p20_data_enable;
  wire p20_not_valid;
  wire p19_enable;
  wire p19_data_enable;
  wire p19_not_valid;
  wire p18_enable;
  wire p18_data_enable;
  wire p18_not_valid;
  wire p17_enable;
  wire p17_data_enable;
  wire p17_not_valid;
  wire p16_enable;
  wire p16_data_enable;
  wire p16_not_valid;
  wire p15_enable;
  wire p15_data_enable;
  wire p15_not_valid;
  wire p14_enable;
  wire p14_data_enable;
  wire p14_not_valid;
  wire p13_enable;
  wire p13_data_enable;
  wire p13_not_valid;
  wire p12_enable;
  wire p12_data_enable;
  wire p12_not_valid;
  wire p11_enable;
  wire p11_data_enable;
  wire p11_not_valid;
  wire p10_enable;
  wire p10_data_enable;
  wire p10_not_valid;
  wire p9_enable;
  wire p9_data_enable;
  wire p9_not_valid;
  wire p8_enable;
  wire p8_data_enable;
  wire p8_not_valid;
  wire p7_enable;
  wire p7_data_enable;
  wire p7_not_valid;
  wire p6_enable;
  wire p6_data_enable;
  wire p6_not_valid;
  wire p5_enable;
  wire p5_data_enable;
  wire p5_not_valid;
  wire p4_enable;
  wire p4_data_enable;
  wire p4_not_valid;
  wire p3_enable;
  wire p3_data_enable;
  wire p3_not_valid;
  wire p2_enable;
  wire p2_data_enable;
  wire p2_not_valid;
  wire p1_enable;
  wire [32:0] r__61;
  wire [31:0] concat_8612;
  wire [31:0] r__92;
  wire [31:0] sub_8364;
  wire [32:0] r__51;
  wire [31:0] concat_8282;
  wire [31:0] r__87;
  wire [31:0] sub_8034;
  wire [32:0] r__41;
  wire [31:0] concat_7952;
  wire [31:0] r__82;
  wire [31:0] sub_7704;
  wire [32:0] r__31;
  wire [31:0] concat_7622;
  wire [31:0] r__77;
  wire [31:0] sub_7374;
  wire [32:0] r__21;
  wire [31:0] concat_7292;
  wire [31:0] r__72;
  wire [31:0] sub_7044;
  wire [32:0] r__11;
  wire [31:0] concat_6962;
  wire [31:0] r__67;
  wire [31:0] sub_6714;
  wire [31:0] concat_6628;
  wire p1_data_enable;
  wire p1_not_valid;
  wire uge_8613;
  wire [31:0] sub_8614;
  wire [32:0] r__59;
  wire [31:0] concat_8530;
  wire [31:0] r__91;
  wire uge_8283;
  wire [31:0] sub_8284;
  wire [32:0] r__49;
  wire [31:0] concat_8200;
  wire [31:0] r__86;
  wire uge_7953;
  wire [31:0] sub_7954;
  wire [32:0] r__39;
  wire [31:0] concat_7870;
  wire [31:0] r__81;
  wire uge_7623;
  wire [31:0] sub_7624;
  wire [32:0] r__29;
  wire [31:0] concat_7540;
  wire [31:0] r__76;
  wire uge_7293;
  wire [31:0] sub_7294;
  wire [32:0] r__19;
  wire [31:0] concat_7210;
  wire [31:0] r__71;
  wire uge_6963;
  wire [31:0] sub_6964;
  wire [32:0] r__9;
  wire [31:0] concat_6880;
  wire [31:0] r__66;
  wire uge_6629;
  wire [31:0] sub_6630;
  wire p0_enable;
  wire p0_all_active_inputs_valid;
  wire [31:0] r__95;
  wire uge_8531;
  wire [31:0] sub_8532;
  wire [32:0] r__57;
  wire [31:0] concat_8450;
  wire [31:0] r__90;
  wire uge_8201;
  wire [31:0] sub_8202;
  wire [32:0] r__47;
  wire [31:0] concat_8120;
  wire [31:0] r__85;
  wire uge_7871;
  wire [31:0] sub_7872;
  wire [32:0] r__37;
  wire [31:0] concat_7790;
  wire [31:0] r__80;
  wire uge_7541;
  wire [31:0] sub_7542;
  wire [32:0] r__27;
  wire [31:0] concat_7460;
  wire [31:0] r__75;
  wire uge_7211;
  wire [31:0] sub_7212;
  wire [32:0] r__17;
  wire [31:0] concat_7130;
  wire [31:0] r__70;
  wire uge_6881;
  wire [31:0] sub_6882;
  wire [32:0] r__7;
  wire [31:0] concat_6800;
  wire [31:0] r__65;
  wire p0_data_enable;
  wire lhs_valid_inv;
  wire rhs_valid_inv;
  wire [31:0] q__32;
  wire [32:0] r__63;
  wire [31:0] r__94;
  wire uge_8451;
  wire [31:0] sub_8452;
  wire [32:0] r__55;
  wire [31:0] concat_8368;
  wire [32:0] r__53;
  wire [31:0] r__89;
  wire uge_8121;
  wire [31:0] sub_8122;
  wire [32:0] r__45;
  wire [31:0] concat_8038;
  wire [32:0] r__43;
  wire [31:0] r__84;
  wire uge_7791;
  wire [31:0] sub_7792;
  wire [32:0] r__35;
  wire [31:0] concat_7708;
  wire [32:0] r__33;
  wire [31:0] r__79;
  wire uge_7461;
  wire [31:0] sub_7462;
  wire [32:0] r__25;
  wire [31:0] concat_7378;
  wire [32:0] r__23;
  wire [31:0] r__74;
  wire uge_7131;
  wire [31:0] sub_7132;
  wire [32:0] r__15;
  wire [31:0] concat_7048;
  wire [32:0] r__13;
  wire [31:0] r__69;
  wire uge_6801;
  wire [31:0] sub_6802;
  wire [32:0] r__5;
  wire [31:0] concat_6718;
  wire [32:0] r__3;
  wire [32:0] bivisor__1;
  wire sign_b;
  wire lhs_valid_load_en;
  wire rhs_valid_load_en;
  wire p30_enable;
  wire p29_enable;
  wire p28_enable;
  wire p27_enable;
  wire p26_enable;
  wire q__32_squeezed_portion_0_width_1;
  wire [30:0] bit_slice_8534;
  wire [31:0] r__93;
  wire uge_8369;
  wire [31:0] sub_8370;
  wire [31:0] concat_8288;
  wire uge_8289;
  wire [30:0] bit_slice_8204;
  wire [31:0] r__88;
  wire uge_8039;
  wire [31:0] sub_8040;
  wire [31:0] concat_7958;
  wire uge_7959;
  wire [30:0] bit_slice_7874;
  wire [31:0] r__83;
  wire uge_7709;
  wire [31:0] sub_7710;
  wire [31:0] concat_7628;
  wire uge_7629;
  wire [30:0] bit_slice_7544;
  wire [31:0] r__78;
  wire uge_7379;
  wire [31:0] sub_7380;
  wire [31:0] concat_7298;
  wire uge_7299;
  wire [30:0] bit_slice_7214;
  wire [31:0] r__73;
  wire uge_7049;
  wire [31:0] sub_7050;
  wire [31:0] concat_6968;
  wire uge_6969;
  wire [30:0] bit_slice_6884;
  wire [31:0] r__68;
  wire uge_6719;
  wire [31:0] sub_6720;
  wire [31:0] concat_6636;
  wire uge_6637;
  wire negated;
  wire sign_a;
  wire bit_slice_6525;
  wire bit_slice_6526;
  wire bit_slice_6527;
  wire bit_slice_6528;
  wire bit_slice_6529;
  wire bit_slice_6530;
  wire bit_slice_6531;
  wire bit_slice_6532;
  wire bit_slice_6533;
  wire bit_slice_6534;
  wire bit_slice_6535;
  wire bit_slice_6536;
  wire bit_slice_6537;
  wire bit_slice_6538;
  wire bit_slice_6539;
  wire bit_slice_6540;
  wire bit_slice_6541;
  wire bit_slice_6542;
  wire bit_slice_6543;
  wire bit_slice_6544;
  wire bit_slice_6545;
  wire bit_slice_6546;
  wire bit_slice_6547;
  wire bit_slice_6548;
  wire bit_slice_6549;
  wire bit_slice_6550;
  wire bit_slice_6551;
  wire bit_slice_6552;
  wire bit_slice_6553;
  wire bit_slice_6554;
  wire bit_slice_6555;
  wire lhs_load_en;
  wire rhs_load_en;
  wire [31:0] signed_div;
  assign result_valid_inv = ~result_valid_reg;
  assign result_valid_load_en = result_ready | result_valid_inv;
  assign result_load_en = p25_valid & result_valid_load_en;
  assign p26_stage_done = p25_valid & result_load_en;
  assign p26_not_valid = ~p25_valid;
  assign p25_enable = p26_stage_done | p26_not_valid;
  assign p25_data_enable = p25_enable & p24_valid;
  assign p25_not_valid = ~p24_valid;
  assign p24_enable = p25_data_enable | p25_not_valid;
  assign p24_data_enable = p24_enable & p23_valid;
  assign p24_not_valid = ~p23_valid;
  assign p23_enable = p24_data_enable | p24_not_valid;
  assign p23_data_enable = p23_enable & p22_valid;
  assign p23_not_valid = ~p22_valid;
  assign p22_enable = p23_data_enable | p23_not_valid;
  assign p22_data_enable = p22_enable & p21_valid;
  assign p22_not_valid = ~p21_valid;
  assign p21_enable = p22_data_enable | p22_not_valid;
  assign p21_data_enable = p21_enable & p20_valid;
  assign p21_not_valid = ~p20_valid;
  assign p20_enable = p21_data_enable | p21_not_valid;
  assign p20_data_enable = p20_enable & p19_valid;
  assign p20_not_valid = ~p19_valid;
  assign p19_enable = p20_data_enable | p20_not_valid;
  assign p19_data_enable = p19_enable & p18_valid;
  assign p19_not_valid = ~p18_valid;
  assign p18_enable = p19_data_enable | p19_not_valid;
  assign p18_data_enable = p18_enable & p17_valid;
  assign p18_not_valid = ~p17_valid;
  assign p17_enable = p18_data_enable | p18_not_valid;
  assign p17_data_enable = p17_enable & p16_valid;
  assign p17_not_valid = ~p16_valid;
  assign p16_enable = p17_data_enable | p17_not_valid;
  assign p16_data_enable = p16_enable & p15_valid;
  assign p16_not_valid = ~p15_valid;
  assign p15_enable = p16_data_enable | p16_not_valid;
  assign p15_data_enable = p15_enable & p14_valid;
  assign p15_not_valid = ~p14_valid;
  assign p14_enable = p15_data_enable | p15_not_valid;
  assign p14_data_enable = p14_enable & p13_valid;
  assign p14_not_valid = ~p13_valid;
  assign p13_enable = p14_data_enable | p14_not_valid;
  assign p13_data_enable = p13_enable & p12_valid;
  assign p13_not_valid = ~p12_valid;
  assign p12_enable = p13_data_enable | p13_not_valid;
  assign p12_data_enable = p12_enable & p11_valid;
  assign p12_not_valid = ~p11_valid;
  assign p11_enable = p12_data_enable | p12_not_valid;
  assign p11_data_enable = p11_enable & p10_valid;
  assign p11_not_valid = ~p10_valid;
  assign p10_enable = p11_data_enable | p11_not_valid;
  assign p10_data_enable = p10_enable & p9_valid;
  assign p10_not_valid = ~p9_valid;
  assign p9_enable = p10_data_enable | p10_not_valid;
  assign p9_data_enable = p9_enable & p8_valid;
  assign p9_not_valid = ~p8_valid;
  assign p8_enable = p9_data_enable | p9_not_valid;
  assign p8_data_enable = p8_enable & p7_valid;
  assign p8_not_valid = ~p7_valid;
  assign p7_enable = p8_data_enable | p8_not_valid;
  assign p7_data_enable = p7_enable & p6_valid;
  assign p7_not_valid = ~p6_valid;
  assign p6_enable = p7_data_enable | p7_not_valid;
  assign p6_data_enable = p6_enable & p5_valid;
  assign p6_not_valid = ~p5_valid;
  assign p5_enable = p6_data_enable | p6_not_valid;
  assign p5_data_enable = p5_enable & p4_valid;
  assign p5_not_valid = ~p4_valid;
  assign p4_enable = p5_data_enable | p5_not_valid;
  assign p4_data_enable = p4_enable & p3_valid;
  assign p4_not_valid = ~p3_valid;
  assign p3_enable = p4_data_enable | p4_not_valid;
  assign p3_data_enable = p3_enable & p2_valid;
  assign p3_not_valid = ~p2_valid;
  assign p2_enable = p3_data_enable | p3_not_valid;
  assign p2_data_enable = p2_enable & p1_valid;
  assign p2_not_valid = ~p1_valid;
  assign p1_enable = p2_data_enable | p2_not_valid;
  assign r__61 = {p24_r__94, p24_bit_slice_6554};
  assign concat_8612 = {p24_bit_slice_8534, p24_bit_slice_6554};
  assign r__92 = p22_uge_8369 ? p22_sub_8370 : p22_concat_8368;
  assign sub_8364 = p21_concat_8288 - p21_b;
  assign r__51 = {p20_r__89, p20_bit_slice_6549};
  assign concat_8282 = {p20_bit_slice_8204, p20_bit_slice_6549};
  assign r__87 = p18_uge_8039 ? p18_sub_8040 : p18_concat_8038;
  assign sub_8034 = p17_concat_7958 - p17_b;
  assign r__41 = {p16_r__84, p16_bit_slice_6544};
  assign concat_7952 = {p16_bit_slice_7874, p16_bit_slice_6544};
  assign r__82 = p14_uge_7709 ? p14_sub_7710 : p14_concat_7708;
  assign sub_7704 = p13_concat_7628 - p13_b;
  assign r__31 = {p12_r__79, p12_bit_slice_6539};
  assign concat_7622 = {p12_bit_slice_7544, p12_bit_slice_6539};
  assign r__77 = p10_uge_7379 ? p10_sub_7380 : p10_concat_7378;
  assign sub_7374 = p9_concat_7298 - p9_b;
  assign r__21 = {p8_r__74, p8_bit_slice_6534};
  assign concat_7292 = {p8_bit_slice_7214, p8_bit_slice_6534};
  assign r__72 = p6_uge_7049 ? p6_sub_7050 : p6_concat_7048;
  assign sub_7044 = p5_concat_6968 - p5_b;
  assign r__11 = {p4_r__69, p4_bit_slice_6529};
  assign concat_6962 = {p4_bit_slice_6884, p4_bit_slice_6529};
  assign r__67 = p2_uge_6719 ? p2_sub_6720 : p2_concat_6718;
  assign sub_6714 = p1_concat_6636 - p1_b;
  assign concat_6628 = {31'h0000_0000, p0_sign_a};
  assign p1_data_enable = p1_enable & p0_valid;
  assign p1_not_valid = ~p0_valid;
  assign uge_8613 = r__61 >= p24_bivisor__1;
  assign sub_8614 = concat_8612 - p24_b;
  assign r__59 = {p23_r__93, p23_bit_slice_6553};
  assign concat_8530 = {p23_r__93[30:0], p23_bit_slice_6553};
  assign r__91 = p21_uge_8289 ? sub_8364 : p21_concat_8288;
  assign uge_8283 = r__51 >= p20_bivisor__1;
  assign sub_8284 = concat_8282 - p20_b;
  assign r__49 = {p19_r__88, p19_bit_slice_6548};
  assign concat_8200 = {p19_r__88[30:0], p19_bit_slice_6548};
  assign r__86 = p17_uge_7959 ? sub_8034 : p17_concat_7958;
  assign uge_7953 = r__41 >= p16_bivisor__1;
  assign sub_7954 = concat_7952 - p16_b;
  assign r__39 = {p15_r__83, p15_bit_slice_6543};
  assign concat_7870 = {p15_r__83[30:0], p15_bit_slice_6543};
  assign r__81 = p13_uge_7629 ? sub_7704 : p13_concat_7628;
  assign uge_7623 = r__31 >= p12_bivisor__1;
  assign sub_7624 = concat_7622 - p12_b;
  assign r__29 = {p11_r__78, p11_bit_slice_6538};
  assign concat_7540 = {p11_r__78[30:0], p11_bit_slice_6538};
  assign r__76 = p9_uge_7299 ? sub_7374 : p9_concat_7298;
  assign uge_7293 = r__21 >= p8_bivisor__1;
  assign sub_7294 = concat_7292 - p8_b;
  assign r__19 = {p7_r__73, p7_bit_slice_6533};
  assign concat_7210 = {p7_r__73[30:0], p7_bit_slice_6533};
  assign r__71 = p5_uge_6969 ? sub_7044 : p5_concat_6968;
  assign uge_6963 = r__11 >= p4_bivisor__1;
  assign sub_6964 = concat_6962 - p4_b;
  assign r__9 = {p3_r__68, p3_bit_slice_6528};
  assign concat_6880 = {p3_r__68[30:0], p3_bit_slice_6528};
  assign r__66 = p1_uge_6637 ? sub_6714 : p1_concat_6636;
  assign uge_6629 = concat_6628 >= p0_b;
  assign sub_6630 = concat_6628 - p0_b;
  assign p0_enable = p1_data_enable | p1_not_valid;
  assign p0_all_active_inputs_valid = lhs_valid_reg & rhs_valid_reg;
  assign r__95 = uge_8613 ? sub_8614 : concat_8612;
  assign uge_8531 = r__59 >= p23_bivisor__1;
  assign sub_8532 = concat_8530 - p23_b;
  assign r__57 = {r__92, p22_bit_slice_6552};
  assign concat_8450 = {r__92[30:0], p22_bit_slice_6552};
  assign r__90 = uge_8283 ? sub_8284 : concat_8282;
  assign uge_8201 = r__49 >= p19_bivisor__1;
  assign sub_8202 = concat_8200 - p19_b;
  assign r__47 = {r__87, p18_bit_slice_6547};
  assign concat_8120 = {r__87[30:0], p18_bit_slice_6547};
  assign r__85 = uge_7953 ? sub_7954 : concat_7952;
  assign uge_7871 = r__39 >= p15_bivisor__1;
  assign sub_7872 = concat_7870 - p15_b;
  assign r__37 = {r__82, p14_bit_slice_6542};
  assign concat_7790 = {r__82[30:0], p14_bit_slice_6542};
  assign r__80 = uge_7623 ? sub_7624 : concat_7622;
  assign uge_7541 = r__29 >= p11_bivisor__1;
  assign sub_7542 = concat_7540 - p11_b;
  assign r__27 = {r__77, p10_bit_slice_6537};
  assign concat_7460 = {r__77[30:0], p10_bit_slice_6537};
  assign r__75 = uge_7293 ? sub_7294 : concat_7292;
  assign uge_7211 = r__19 >= p7_bivisor__1;
  assign sub_7212 = concat_7210 - p7_b;
  assign r__17 = {r__72, p6_bit_slice_6532};
  assign concat_7130 = {r__72[30:0], p6_bit_slice_6532};
  assign r__70 = uge_6963 ? sub_6964 : concat_6962;
  assign uge_6881 = r__9 >= p3_bivisor__1;
  assign sub_6882 = concat_6880 - p3_b;
  assign r__7 = {r__67, p2_bit_slice_6527};
  assign concat_6800 = {r__67[30:0], p2_bit_slice_6527};
  assign r__65 = uge_6629 ? sub_6630 : concat_6628;
  assign p0_data_enable = p0_enable & p0_all_active_inputs_valid;
  assign lhs_valid_inv = ~lhs_valid_reg;
  assign rhs_valid_inv = ~rhs_valid_reg;
  assign q__32 = {p25_uge_6629, p25_uge_6637, p25_uge_6719, p25_uge_6801, p25_uge_6881, p25_uge_6963, p25_uge_6969, p25_uge_7049, p25_uge_7131, p25_uge_7211, p25_uge_7293, p25_uge_7299, p25_uge_7379, p25_uge_7461, p25_uge_7541, p25_uge_7623, p25_uge_7629, p25_uge_7709, p25_uge_7791, p25_uge_7871, p25_uge_7953, p25_uge_7959, p25_uge_8039, p25_uge_8121, p25_uge_8201, p25_uge_8283, p25_uge_8289, p25_uge_8369, p25_uge_8451, p25_uge_8531, p25_uge_8613, p25_q__32_squeezed_portion_0_width_1};
  assign r__63 = {r__95, p24_bit_slice_6555};
  assign r__94 = uge_8531 ? sub_8532 : concat_8530;
  assign uge_8451 = r__57 >= p22_bivisor__1;
  assign sub_8452 = concat_8450 - p22_b;
  assign r__55 = {r__91, p21_bit_slice_6551};
  assign concat_8368 = {r__91[30:0], p21_bit_slice_6551};
  assign r__53 = {r__90, p20_bit_slice_6550};
  assign r__89 = uge_8201 ? sub_8202 : concat_8200;
  assign uge_8121 = r__47 >= p18_bivisor__1;
  assign sub_8122 = concat_8120 - p18_b;
  assign r__45 = {r__86, p17_bit_slice_6546};
  assign concat_8038 = {r__86[30:0], p17_bit_slice_6546};
  assign r__43 = {r__85, p16_bit_slice_6545};
  assign r__84 = uge_7871 ? sub_7872 : concat_7870;
  assign uge_7791 = r__37 >= p14_bivisor__1;
  assign sub_7792 = concat_7790 - p14_b;
  assign r__35 = {r__81, p13_bit_slice_6541};
  assign concat_7708 = {r__81[30:0], p13_bit_slice_6541};
  assign r__33 = {r__80, p12_bit_slice_6540};
  assign r__79 = uge_7541 ? sub_7542 : concat_7540;
  assign uge_7461 = r__27 >= p10_bivisor__1;
  assign sub_7462 = concat_7460 - p10_b;
  assign r__25 = {r__76, p9_bit_slice_6536};
  assign concat_7378 = {r__76[30:0], p9_bit_slice_6536};
  assign r__23 = {r__75, p8_bit_slice_6535};
  assign r__74 = uge_7211 ? sub_7212 : concat_7210;
  assign uge_7131 = r__17 >= p6_bivisor__1;
  assign sub_7132 = concat_7130 - p6_b;
  assign r__15 = {r__71, p5_bit_slice_6531};
  assign concat_7048 = {r__71[30:0], p5_bit_slice_6531};
  assign r__13 = {r__70, p4_bit_slice_6530};
  assign r__69 = uge_6881 ? sub_6882 : concat_6880;
  assign uge_6801 = r__7 >= p2_bivisor__1;
  assign sub_6802 = concat_6800 - p2_b;
  assign r__5 = {r__66, p1_bit_slice_6526};
  assign concat_6718 = {r__66[30:0], p1_bit_slice_6526};
  assign r__3 = {r__65, p0_bit_slice_6525};
  assign bivisor__1 = {1'h0, p0_b};
  assign sign_b = p0_b[31];
  assign lhs_valid_load_en = p0_data_enable | lhs_valid_inv;
  assign rhs_valid_load_en = p0_data_enable | rhs_valid_inv;
  assign p30_enable = 1'h1;
  assign p29_enable = 1'h1;
  assign p28_enable = 1'h1;
  assign p27_enable = 1'h1;
  assign p26_enable = 1'h1;
  assign q__32_squeezed_portion_0_width_1 = r__63 >= p24_bivisor__1;
  assign bit_slice_8534 = r__94[30:0];
  assign r__93 = uge_8451 ? sub_8452 : concat_8450;
  assign uge_8369 = r__55 >= p21_bivisor__1;
  assign sub_8370 = concat_8368 - p21_b;
  assign concat_8288 = {r__90[30:0], p20_bit_slice_6550};
  assign uge_8289 = r__53 >= p20_bivisor__1;
  assign bit_slice_8204 = r__89[30:0];
  assign r__88 = uge_8121 ? sub_8122 : concat_8120;
  assign uge_8039 = r__45 >= p17_bivisor__1;
  assign sub_8040 = concat_8038 - p17_b;
  assign concat_7958 = {r__85[30:0], p16_bit_slice_6545};
  assign uge_7959 = r__43 >= p16_bivisor__1;
  assign bit_slice_7874 = r__84[30:0];
  assign r__83 = uge_7791 ? sub_7792 : concat_7790;
  assign uge_7709 = r__35 >= p13_bivisor__1;
  assign sub_7710 = concat_7708 - p13_b;
  assign concat_7628 = {r__80[30:0], p12_bit_slice_6540};
  assign uge_7629 = r__33 >= p12_bivisor__1;
  assign bit_slice_7544 = r__79[30:0];
  assign r__78 = uge_7461 ? sub_7462 : concat_7460;
  assign uge_7379 = r__25 >= p9_bivisor__1;
  assign sub_7380 = concat_7378 - p9_b;
  assign concat_7298 = {r__75[30:0], p8_bit_slice_6535};
  assign uge_7299 = r__23 >= p8_bivisor__1;
  assign bit_slice_7214 = r__74[30:0];
  assign r__73 = uge_7131 ? sub_7132 : concat_7130;
  assign uge_7049 = r__15 >= p5_bivisor__1;
  assign sub_7050 = concat_7048 - p5_b;
  assign concat_6968 = {r__70[30:0], p4_bit_slice_6530};
  assign uge_6969 = r__13 >= p4_bivisor__1;
  assign bit_slice_6884 = r__69[30:0];
  assign r__68 = uge_6801 ? sub_6802 : concat_6800;
  assign uge_6719 = r__5 >= p1_bivisor__1;
  assign sub_6720 = concat_6718 - p1_b;
  assign concat_6636 = {r__65[30:0], p0_bit_slice_6525};
  assign uge_6637 = r__3 >= bivisor__1;
  assign negated = p0_sign_a ^ sign_b;
  assign sign_a = lhs_reg[31];
  assign bit_slice_6525 = lhs_reg[30];
  assign bit_slice_6526 = lhs_reg[29];
  assign bit_slice_6527 = lhs_reg[28];
  assign bit_slice_6528 = lhs_reg[27];
  assign bit_slice_6529 = lhs_reg[26];
  assign bit_slice_6530 = lhs_reg[25];
  assign bit_slice_6531 = lhs_reg[24];
  assign bit_slice_6532 = lhs_reg[23];
  assign bit_slice_6533 = lhs_reg[22];
  assign bit_slice_6534 = lhs_reg[21];
  assign bit_slice_6535 = lhs_reg[20];
  assign bit_slice_6536 = lhs_reg[19];
  assign bit_slice_6537 = lhs_reg[18];
  assign bit_slice_6538 = lhs_reg[17];
  assign bit_slice_6539 = lhs_reg[16];
  assign bit_slice_6540 = lhs_reg[15];
  assign bit_slice_6541 = lhs_reg[14];
  assign bit_slice_6542 = lhs_reg[13];
  assign bit_slice_6543 = lhs_reg[12];
  assign bit_slice_6544 = lhs_reg[11];
  assign bit_slice_6545 = lhs_reg[10];
  assign bit_slice_6546 = lhs_reg[9];
  assign bit_slice_6547 = lhs_reg[8];
  assign bit_slice_6548 = lhs_reg[7];
  assign bit_slice_6549 = lhs_reg[6];
  assign bit_slice_6550 = lhs_reg[5];
  assign bit_slice_6551 = lhs_reg[4];
  assign bit_slice_6552 = lhs_reg[3];
  assign bit_slice_6553 = lhs_reg[2];
  assign bit_slice_6554 = lhs_reg[1];
  assign bit_slice_6555 = lhs_reg[0];
  assign lhs_load_en = lhs_valid & lhs_valid_load_en;
  assign rhs_load_en = rhs_valid & rhs_valid_load_en;
  assign signed_div = p25_negated ? -q__32 : q__32;
  always @ (posedge clk) begin
    if (rst) begin
      p0_sign_a <= 1'h0;
      p0_b <= 32'h0000_0000;
      p0_bit_slice_6525 <= 1'h0;
      p0_bit_slice_6526 <= 1'h0;
      p0_bit_slice_6527 <= 1'h0;
      p0_bit_slice_6528 <= 1'h0;
      p0_bit_slice_6529 <= 1'h0;
      p0_bit_slice_6530 <= 1'h0;
      p0_bit_slice_6531 <= 1'h0;
      p0_bit_slice_6532 <= 1'h0;
      p0_bit_slice_6533 <= 1'h0;
      p0_bit_slice_6534 <= 1'h0;
      p0_bit_slice_6535 <= 1'h0;
      p0_bit_slice_6536 <= 1'h0;
      p0_bit_slice_6537 <= 1'h0;
      p0_bit_slice_6538 <= 1'h0;
      p0_bit_slice_6539 <= 1'h0;
      p0_bit_slice_6540 <= 1'h0;
      p0_bit_slice_6541 <= 1'h0;
      p0_bit_slice_6542 <= 1'h0;
      p0_bit_slice_6543 <= 1'h0;
      p0_bit_slice_6544 <= 1'h0;
      p0_bit_slice_6545 <= 1'h0;
      p0_bit_slice_6546 <= 1'h0;
      p0_bit_slice_6547 <= 1'h0;
      p0_bit_slice_6548 <= 1'h0;
      p0_bit_slice_6549 <= 1'h0;
      p0_bit_slice_6550 <= 1'h0;
      p0_bit_slice_6551 <= 1'h0;
      p0_bit_slice_6552 <= 1'h0;
      p0_bit_slice_6553 <= 1'h0;
      p0_bit_slice_6554 <= 1'h0;
      p0_bit_slice_6555 <= 1'h0;
      p1_b <= 32'h0000_0000;
      p1_uge_6629 <= 1'h0;
      p1_bivisor__1 <= 33'h0_0000_0000;
      p1_concat_6636 <= 32'h0000_0000;
      p1_uge_6637 <= 1'h0;
      p1_bit_slice_6526 <= 1'h0;
      p1_bit_slice_6527 <= 1'h0;
      p1_bit_slice_6528 <= 1'h0;
      p1_bit_slice_6529 <= 1'h0;
      p1_bit_slice_6530 <= 1'h0;
      p1_bit_slice_6531 <= 1'h0;
      p1_bit_slice_6532 <= 1'h0;
      p1_bit_slice_6533 <= 1'h0;
      p1_bit_slice_6534 <= 1'h0;
      p1_bit_slice_6535 <= 1'h0;
      p1_bit_slice_6536 <= 1'h0;
      p1_bit_slice_6537 <= 1'h0;
      p1_bit_slice_6538 <= 1'h0;
      p1_bit_slice_6539 <= 1'h0;
      p1_bit_slice_6540 <= 1'h0;
      p1_bit_slice_6541 <= 1'h0;
      p1_bit_slice_6542 <= 1'h0;
      p1_bit_slice_6543 <= 1'h0;
      p1_bit_slice_6544 <= 1'h0;
      p1_bit_slice_6545 <= 1'h0;
      p1_bit_slice_6546 <= 1'h0;
      p1_bit_slice_6547 <= 1'h0;
      p1_bit_slice_6548 <= 1'h0;
      p1_bit_slice_6549 <= 1'h0;
      p1_bit_slice_6550 <= 1'h0;
      p1_bit_slice_6551 <= 1'h0;
      p1_bit_slice_6552 <= 1'h0;
      p1_bit_slice_6553 <= 1'h0;
      p1_bit_slice_6554 <= 1'h0;
      p1_bit_slice_6555 <= 1'h0;
      p1_negated <= 1'h0;
      p2_b <= 32'h0000_0000;
      p2_uge_6629 <= 1'h0;
      p2_bivisor__1 <= 33'h0_0000_0000;
      p2_uge_6637 <= 1'h0;
      p2_concat_6718 <= 32'h0000_0000;
      p2_uge_6719 <= 1'h0;
      p2_sub_6720 <= 32'h0000_0000;
      p2_bit_slice_6527 <= 1'h0;
      p2_bit_slice_6528 <= 1'h0;
      p2_bit_slice_6529 <= 1'h0;
      p2_bit_slice_6530 <= 1'h0;
      p2_bit_slice_6531 <= 1'h0;
      p2_bit_slice_6532 <= 1'h0;
      p2_bit_slice_6533 <= 1'h0;
      p2_bit_slice_6534 <= 1'h0;
      p2_bit_slice_6535 <= 1'h0;
      p2_bit_slice_6536 <= 1'h0;
      p2_bit_slice_6537 <= 1'h0;
      p2_bit_slice_6538 <= 1'h0;
      p2_bit_slice_6539 <= 1'h0;
      p2_bit_slice_6540 <= 1'h0;
      p2_bit_slice_6541 <= 1'h0;
      p2_bit_slice_6542 <= 1'h0;
      p2_bit_slice_6543 <= 1'h0;
      p2_bit_slice_6544 <= 1'h0;
      p2_bit_slice_6545 <= 1'h0;
      p2_bit_slice_6546 <= 1'h0;
      p2_bit_slice_6547 <= 1'h0;
      p2_bit_slice_6548 <= 1'h0;
      p2_bit_slice_6549 <= 1'h0;
      p2_bit_slice_6550 <= 1'h0;
      p2_bit_slice_6551 <= 1'h0;
      p2_bit_slice_6552 <= 1'h0;
      p2_bit_slice_6553 <= 1'h0;
      p2_bit_slice_6554 <= 1'h0;
      p2_bit_slice_6555 <= 1'h0;
      p2_negated <= 1'h0;
      p3_b <= 32'h0000_0000;
      p3_uge_6629 <= 1'h0;
      p3_bivisor__1 <= 33'h0_0000_0000;
      p3_uge_6637 <= 1'h0;
      p3_uge_6719 <= 1'h0;
      p3_uge_6801 <= 1'h0;
      p3_r__68 <= 32'h0000_0000;
      p3_bit_slice_6528 <= 1'h0;
      p3_bit_slice_6529 <= 1'h0;
      p3_bit_slice_6530 <= 1'h0;
      p3_bit_slice_6531 <= 1'h0;
      p3_bit_slice_6532 <= 1'h0;
      p3_bit_slice_6533 <= 1'h0;
      p3_bit_slice_6534 <= 1'h0;
      p3_bit_slice_6535 <= 1'h0;
      p3_bit_slice_6536 <= 1'h0;
      p3_bit_slice_6537 <= 1'h0;
      p3_bit_slice_6538 <= 1'h0;
      p3_bit_slice_6539 <= 1'h0;
      p3_bit_slice_6540 <= 1'h0;
      p3_bit_slice_6541 <= 1'h0;
      p3_bit_slice_6542 <= 1'h0;
      p3_bit_slice_6543 <= 1'h0;
      p3_bit_slice_6544 <= 1'h0;
      p3_bit_slice_6545 <= 1'h0;
      p3_bit_slice_6546 <= 1'h0;
      p3_bit_slice_6547 <= 1'h0;
      p3_bit_slice_6548 <= 1'h0;
      p3_bit_slice_6549 <= 1'h0;
      p3_bit_slice_6550 <= 1'h0;
      p3_bit_slice_6551 <= 1'h0;
      p3_bit_slice_6552 <= 1'h0;
      p3_bit_slice_6553 <= 1'h0;
      p3_bit_slice_6554 <= 1'h0;
      p3_bit_slice_6555 <= 1'h0;
      p3_negated <= 1'h0;
      p4_b <= 32'h0000_0000;
      p4_uge_6629 <= 1'h0;
      p4_bivisor__1 <= 33'h0_0000_0000;
      p4_uge_6637 <= 1'h0;
      p4_uge_6719 <= 1'h0;
      p4_uge_6801 <= 1'h0;
      p4_uge_6881 <= 1'h0;
      p4_r__69 <= 32'h0000_0000;
      p4_bit_slice_6529 <= 1'h0;
      p4_bit_slice_6884 <= 31'h0000_0000;
      p4_bit_slice_6530 <= 1'h0;
      p4_bit_slice_6531 <= 1'h0;
      p4_bit_slice_6532 <= 1'h0;
      p4_bit_slice_6533 <= 1'h0;
      p4_bit_slice_6534 <= 1'h0;
      p4_bit_slice_6535 <= 1'h0;
      p4_bit_slice_6536 <= 1'h0;
      p4_bit_slice_6537 <= 1'h0;
      p4_bit_slice_6538 <= 1'h0;
      p4_bit_slice_6539 <= 1'h0;
      p4_bit_slice_6540 <= 1'h0;
      p4_bit_slice_6541 <= 1'h0;
      p4_bit_slice_6542 <= 1'h0;
      p4_bit_slice_6543 <= 1'h0;
      p4_bit_slice_6544 <= 1'h0;
      p4_bit_slice_6545 <= 1'h0;
      p4_bit_slice_6546 <= 1'h0;
      p4_bit_slice_6547 <= 1'h0;
      p4_bit_slice_6548 <= 1'h0;
      p4_bit_slice_6549 <= 1'h0;
      p4_bit_slice_6550 <= 1'h0;
      p4_bit_slice_6551 <= 1'h0;
      p4_bit_slice_6552 <= 1'h0;
      p4_bit_slice_6553 <= 1'h0;
      p4_bit_slice_6554 <= 1'h0;
      p4_bit_slice_6555 <= 1'h0;
      p4_negated <= 1'h0;
      p5_b <= 32'h0000_0000;
      p5_uge_6629 <= 1'h0;
      p5_bivisor__1 <= 33'h0_0000_0000;
      p5_uge_6637 <= 1'h0;
      p5_uge_6719 <= 1'h0;
      p5_uge_6801 <= 1'h0;
      p5_uge_6881 <= 1'h0;
      p5_uge_6963 <= 1'h0;
      p5_concat_6968 <= 32'h0000_0000;
      p5_uge_6969 <= 1'h0;
      p5_bit_slice_6531 <= 1'h0;
      p5_bit_slice_6532 <= 1'h0;
      p5_bit_slice_6533 <= 1'h0;
      p5_bit_slice_6534 <= 1'h0;
      p5_bit_slice_6535 <= 1'h0;
      p5_bit_slice_6536 <= 1'h0;
      p5_bit_slice_6537 <= 1'h0;
      p5_bit_slice_6538 <= 1'h0;
      p5_bit_slice_6539 <= 1'h0;
      p5_bit_slice_6540 <= 1'h0;
      p5_bit_slice_6541 <= 1'h0;
      p5_bit_slice_6542 <= 1'h0;
      p5_bit_slice_6543 <= 1'h0;
      p5_bit_slice_6544 <= 1'h0;
      p5_bit_slice_6545 <= 1'h0;
      p5_bit_slice_6546 <= 1'h0;
      p5_bit_slice_6547 <= 1'h0;
      p5_bit_slice_6548 <= 1'h0;
      p5_bit_slice_6549 <= 1'h0;
      p5_bit_slice_6550 <= 1'h0;
      p5_bit_slice_6551 <= 1'h0;
      p5_bit_slice_6552 <= 1'h0;
      p5_bit_slice_6553 <= 1'h0;
      p5_bit_slice_6554 <= 1'h0;
      p5_bit_slice_6555 <= 1'h0;
      p5_negated <= 1'h0;
      p6_b <= 32'h0000_0000;
      p6_uge_6629 <= 1'h0;
      p6_bivisor__1 <= 33'h0_0000_0000;
      p6_uge_6637 <= 1'h0;
      p6_uge_6719 <= 1'h0;
      p6_uge_6801 <= 1'h0;
      p6_uge_6881 <= 1'h0;
      p6_uge_6963 <= 1'h0;
      p6_uge_6969 <= 1'h0;
      p6_concat_7048 <= 32'h0000_0000;
      p6_uge_7049 <= 1'h0;
      p6_sub_7050 <= 32'h0000_0000;
      p6_bit_slice_6532 <= 1'h0;
      p6_bit_slice_6533 <= 1'h0;
      p6_bit_slice_6534 <= 1'h0;
      p6_bit_slice_6535 <= 1'h0;
      p6_bit_slice_6536 <= 1'h0;
      p6_bit_slice_6537 <= 1'h0;
      p6_bit_slice_6538 <= 1'h0;
      p6_bit_slice_6539 <= 1'h0;
      p6_bit_slice_6540 <= 1'h0;
      p6_bit_slice_6541 <= 1'h0;
      p6_bit_slice_6542 <= 1'h0;
      p6_bit_slice_6543 <= 1'h0;
      p6_bit_slice_6544 <= 1'h0;
      p6_bit_slice_6545 <= 1'h0;
      p6_bit_slice_6546 <= 1'h0;
      p6_bit_slice_6547 <= 1'h0;
      p6_bit_slice_6548 <= 1'h0;
      p6_bit_slice_6549 <= 1'h0;
      p6_bit_slice_6550 <= 1'h0;
      p6_bit_slice_6551 <= 1'h0;
      p6_bit_slice_6552 <= 1'h0;
      p6_bit_slice_6553 <= 1'h0;
      p6_bit_slice_6554 <= 1'h0;
      p6_bit_slice_6555 <= 1'h0;
      p6_negated <= 1'h0;
      p7_b <= 32'h0000_0000;
      p7_uge_6629 <= 1'h0;
      p7_bivisor__1 <= 33'h0_0000_0000;
      p7_uge_6637 <= 1'h0;
      p7_uge_6719 <= 1'h0;
      p7_uge_6801 <= 1'h0;
      p7_uge_6881 <= 1'h0;
      p7_uge_6963 <= 1'h0;
      p7_uge_6969 <= 1'h0;
      p7_uge_7049 <= 1'h0;
      p7_uge_7131 <= 1'h0;
      p7_r__73 <= 32'h0000_0000;
      p7_bit_slice_6533 <= 1'h0;
      p7_bit_slice_6534 <= 1'h0;
      p7_bit_slice_6535 <= 1'h0;
      p7_bit_slice_6536 <= 1'h0;
      p7_bit_slice_6537 <= 1'h0;
      p7_bit_slice_6538 <= 1'h0;
      p7_bit_slice_6539 <= 1'h0;
      p7_bit_slice_6540 <= 1'h0;
      p7_bit_slice_6541 <= 1'h0;
      p7_bit_slice_6542 <= 1'h0;
      p7_bit_slice_6543 <= 1'h0;
      p7_bit_slice_6544 <= 1'h0;
      p7_bit_slice_6545 <= 1'h0;
      p7_bit_slice_6546 <= 1'h0;
      p7_bit_slice_6547 <= 1'h0;
      p7_bit_slice_6548 <= 1'h0;
      p7_bit_slice_6549 <= 1'h0;
      p7_bit_slice_6550 <= 1'h0;
      p7_bit_slice_6551 <= 1'h0;
      p7_bit_slice_6552 <= 1'h0;
      p7_bit_slice_6553 <= 1'h0;
      p7_bit_slice_6554 <= 1'h0;
      p7_bit_slice_6555 <= 1'h0;
      p7_negated <= 1'h0;
      p8_b <= 32'h0000_0000;
      p8_uge_6629 <= 1'h0;
      p8_bivisor__1 <= 33'h0_0000_0000;
      p8_uge_6637 <= 1'h0;
      p8_uge_6719 <= 1'h0;
      p8_uge_6801 <= 1'h0;
      p8_uge_6881 <= 1'h0;
      p8_uge_6963 <= 1'h0;
      p8_uge_6969 <= 1'h0;
      p8_uge_7049 <= 1'h0;
      p8_uge_7131 <= 1'h0;
      p8_uge_7211 <= 1'h0;
      p8_r__74 <= 32'h0000_0000;
      p8_bit_slice_6534 <= 1'h0;
      p8_bit_slice_7214 <= 31'h0000_0000;
      p8_bit_slice_6535 <= 1'h0;
      p8_bit_slice_6536 <= 1'h0;
      p8_bit_slice_6537 <= 1'h0;
      p8_bit_slice_6538 <= 1'h0;
      p8_bit_slice_6539 <= 1'h0;
      p8_bit_slice_6540 <= 1'h0;
      p8_bit_slice_6541 <= 1'h0;
      p8_bit_slice_6542 <= 1'h0;
      p8_bit_slice_6543 <= 1'h0;
      p8_bit_slice_6544 <= 1'h0;
      p8_bit_slice_6545 <= 1'h0;
      p8_bit_slice_6546 <= 1'h0;
      p8_bit_slice_6547 <= 1'h0;
      p8_bit_slice_6548 <= 1'h0;
      p8_bit_slice_6549 <= 1'h0;
      p8_bit_slice_6550 <= 1'h0;
      p8_bit_slice_6551 <= 1'h0;
      p8_bit_slice_6552 <= 1'h0;
      p8_bit_slice_6553 <= 1'h0;
      p8_bit_slice_6554 <= 1'h0;
      p8_bit_slice_6555 <= 1'h0;
      p8_negated <= 1'h0;
      p9_b <= 32'h0000_0000;
      p9_uge_6629 <= 1'h0;
      p9_bivisor__1 <= 33'h0_0000_0000;
      p9_uge_6637 <= 1'h0;
      p9_uge_6719 <= 1'h0;
      p9_uge_6801 <= 1'h0;
      p9_uge_6881 <= 1'h0;
      p9_uge_6963 <= 1'h0;
      p9_uge_6969 <= 1'h0;
      p9_uge_7049 <= 1'h0;
      p9_uge_7131 <= 1'h0;
      p9_uge_7211 <= 1'h0;
      p9_uge_7293 <= 1'h0;
      p9_concat_7298 <= 32'h0000_0000;
      p9_uge_7299 <= 1'h0;
      p9_bit_slice_6536 <= 1'h0;
      p9_bit_slice_6537 <= 1'h0;
      p9_bit_slice_6538 <= 1'h0;
      p9_bit_slice_6539 <= 1'h0;
      p9_bit_slice_6540 <= 1'h0;
      p9_bit_slice_6541 <= 1'h0;
      p9_bit_slice_6542 <= 1'h0;
      p9_bit_slice_6543 <= 1'h0;
      p9_bit_slice_6544 <= 1'h0;
      p9_bit_slice_6545 <= 1'h0;
      p9_bit_slice_6546 <= 1'h0;
      p9_bit_slice_6547 <= 1'h0;
      p9_bit_slice_6548 <= 1'h0;
      p9_bit_slice_6549 <= 1'h0;
      p9_bit_slice_6550 <= 1'h0;
      p9_bit_slice_6551 <= 1'h0;
      p9_bit_slice_6552 <= 1'h0;
      p9_bit_slice_6553 <= 1'h0;
      p9_bit_slice_6554 <= 1'h0;
      p9_bit_slice_6555 <= 1'h0;
      p9_negated <= 1'h0;
      p10_b <= 32'h0000_0000;
      p10_uge_6629 <= 1'h0;
      p10_bivisor__1 <= 33'h0_0000_0000;
      p10_uge_6637 <= 1'h0;
      p10_uge_6719 <= 1'h0;
      p10_uge_6801 <= 1'h0;
      p10_uge_6881 <= 1'h0;
      p10_uge_6963 <= 1'h0;
      p10_uge_6969 <= 1'h0;
      p10_uge_7049 <= 1'h0;
      p10_uge_7131 <= 1'h0;
      p10_uge_7211 <= 1'h0;
      p10_uge_7293 <= 1'h0;
      p10_uge_7299 <= 1'h0;
      p10_concat_7378 <= 32'h0000_0000;
      p10_uge_7379 <= 1'h0;
      p10_sub_7380 <= 32'h0000_0000;
      p10_bit_slice_6537 <= 1'h0;
      p10_bit_slice_6538 <= 1'h0;
      p10_bit_slice_6539 <= 1'h0;
      p10_bit_slice_6540 <= 1'h0;
      p10_bit_slice_6541 <= 1'h0;
      p10_bit_slice_6542 <= 1'h0;
      p10_bit_slice_6543 <= 1'h0;
      p10_bit_slice_6544 <= 1'h0;
      p10_bit_slice_6545 <= 1'h0;
      p10_bit_slice_6546 <= 1'h0;
      p10_bit_slice_6547 <= 1'h0;
      p10_bit_slice_6548 <= 1'h0;
      p10_bit_slice_6549 <= 1'h0;
      p10_bit_slice_6550 <= 1'h0;
      p10_bit_slice_6551 <= 1'h0;
      p10_bit_slice_6552 <= 1'h0;
      p10_bit_slice_6553 <= 1'h0;
      p10_bit_slice_6554 <= 1'h0;
      p10_bit_slice_6555 <= 1'h0;
      p10_negated <= 1'h0;
      p11_b <= 32'h0000_0000;
      p11_uge_6629 <= 1'h0;
      p11_bivisor__1 <= 33'h0_0000_0000;
      p11_uge_6637 <= 1'h0;
      p11_uge_6719 <= 1'h0;
      p11_uge_6801 <= 1'h0;
      p11_uge_6881 <= 1'h0;
      p11_uge_6963 <= 1'h0;
      p11_uge_6969 <= 1'h0;
      p11_uge_7049 <= 1'h0;
      p11_uge_7131 <= 1'h0;
      p11_uge_7211 <= 1'h0;
      p11_uge_7293 <= 1'h0;
      p11_uge_7299 <= 1'h0;
      p11_uge_7379 <= 1'h0;
      p11_uge_7461 <= 1'h0;
      p11_r__78 <= 32'h0000_0000;
      p11_bit_slice_6538 <= 1'h0;
      p11_bit_slice_6539 <= 1'h0;
      p11_bit_slice_6540 <= 1'h0;
      p11_bit_slice_6541 <= 1'h0;
      p11_bit_slice_6542 <= 1'h0;
      p11_bit_slice_6543 <= 1'h0;
      p11_bit_slice_6544 <= 1'h0;
      p11_bit_slice_6545 <= 1'h0;
      p11_bit_slice_6546 <= 1'h0;
      p11_bit_slice_6547 <= 1'h0;
      p11_bit_slice_6548 <= 1'h0;
      p11_bit_slice_6549 <= 1'h0;
      p11_bit_slice_6550 <= 1'h0;
      p11_bit_slice_6551 <= 1'h0;
      p11_bit_slice_6552 <= 1'h0;
      p11_bit_slice_6553 <= 1'h0;
      p11_bit_slice_6554 <= 1'h0;
      p11_bit_slice_6555 <= 1'h0;
      p11_negated <= 1'h0;
      p12_b <= 32'h0000_0000;
      p12_uge_6629 <= 1'h0;
      p12_bivisor__1 <= 33'h0_0000_0000;
      p12_uge_6637 <= 1'h0;
      p12_uge_6719 <= 1'h0;
      p12_uge_6801 <= 1'h0;
      p12_uge_6881 <= 1'h0;
      p12_uge_6963 <= 1'h0;
      p12_uge_6969 <= 1'h0;
      p12_uge_7049 <= 1'h0;
      p12_uge_7131 <= 1'h0;
      p12_uge_7211 <= 1'h0;
      p12_uge_7293 <= 1'h0;
      p12_uge_7299 <= 1'h0;
      p12_uge_7379 <= 1'h0;
      p12_uge_7461 <= 1'h0;
      p12_uge_7541 <= 1'h0;
      p12_r__79 <= 32'h0000_0000;
      p12_bit_slice_6539 <= 1'h0;
      p12_bit_slice_7544 <= 31'h0000_0000;
      p12_bit_slice_6540 <= 1'h0;
      p12_bit_slice_6541 <= 1'h0;
      p12_bit_slice_6542 <= 1'h0;
      p12_bit_slice_6543 <= 1'h0;
      p12_bit_slice_6544 <= 1'h0;
      p12_bit_slice_6545 <= 1'h0;
      p12_bit_slice_6546 <= 1'h0;
      p12_bit_slice_6547 <= 1'h0;
      p12_bit_slice_6548 <= 1'h0;
      p12_bit_slice_6549 <= 1'h0;
      p12_bit_slice_6550 <= 1'h0;
      p12_bit_slice_6551 <= 1'h0;
      p12_bit_slice_6552 <= 1'h0;
      p12_bit_slice_6553 <= 1'h0;
      p12_bit_slice_6554 <= 1'h0;
      p12_bit_slice_6555 <= 1'h0;
      p12_negated <= 1'h0;
      p13_b <= 32'h0000_0000;
      p13_uge_6629 <= 1'h0;
      p13_bivisor__1 <= 33'h0_0000_0000;
      p13_uge_6637 <= 1'h0;
      p13_uge_6719 <= 1'h0;
      p13_uge_6801 <= 1'h0;
      p13_uge_6881 <= 1'h0;
      p13_uge_6963 <= 1'h0;
      p13_uge_6969 <= 1'h0;
      p13_uge_7049 <= 1'h0;
      p13_uge_7131 <= 1'h0;
      p13_uge_7211 <= 1'h0;
      p13_uge_7293 <= 1'h0;
      p13_uge_7299 <= 1'h0;
      p13_uge_7379 <= 1'h0;
      p13_uge_7461 <= 1'h0;
      p13_uge_7541 <= 1'h0;
      p13_uge_7623 <= 1'h0;
      p13_concat_7628 <= 32'h0000_0000;
      p13_uge_7629 <= 1'h0;
      p13_bit_slice_6541 <= 1'h0;
      p13_bit_slice_6542 <= 1'h0;
      p13_bit_slice_6543 <= 1'h0;
      p13_bit_slice_6544 <= 1'h0;
      p13_bit_slice_6545 <= 1'h0;
      p13_bit_slice_6546 <= 1'h0;
      p13_bit_slice_6547 <= 1'h0;
      p13_bit_slice_6548 <= 1'h0;
      p13_bit_slice_6549 <= 1'h0;
      p13_bit_slice_6550 <= 1'h0;
      p13_bit_slice_6551 <= 1'h0;
      p13_bit_slice_6552 <= 1'h0;
      p13_bit_slice_6553 <= 1'h0;
      p13_bit_slice_6554 <= 1'h0;
      p13_bit_slice_6555 <= 1'h0;
      p13_negated <= 1'h0;
      p14_b <= 32'h0000_0000;
      p14_uge_6629 <= 1'h0;
      p14_bivisor__1 <= 33'h0_0000_0000;
      p14_uge_6637 <= 1'h0;
      p14_uge_6719 <= 1'h0;
      p14_uge_6801 <= 1'h0;
      p14_uge_6881 <= 1'h0;
      p14_uge_6963 <= 1'h0;
      p14_uge_6969 <= 1'h0;
      p14_uge_7049 <= 1'h0;
      p14_uge_7131 <= 1'h0;
      p14_uge_7211 <= 1'h0;
      p14_uge_7293 <= 1'h0;
      p14_uge_7299 <= 1'h0;
      p14_uge_7379 <= 1'h0;
      p14_uge_7461 <= 1'h0;
      p14_uge_7541 <= 1'h0;
      p14_uge_7623 <= 1'h0;
      p14_uge_7629 <= 1'h0;
      p14_concat_7708 <= 32'h0000_0000;
      p14_uge_7709 <= 1'h0;
      p14_sub_7710 <= 32'h0000_0000;
      p14_bit_slice_6542 <= 1'h0;
      p14_bit_slice_6543 <= 1'h0;
      p14_bit_slice_6544 <= 1'h0;
      p14_bit_slice_6545 <= 1'h0;
      p14_bit_slice_6546 <= 1'h0;
      p14_bit_slice_6547 <= 1'h0;
      p14_bit_slice_6548 <= 1'h0;
      p14_bit_slice_6549 <= 1'h0;
      p14_bit_slice_6550 <= 1'h0;
      p14_bit_slice_6551 <= 1'h0;
      p14_bit_slice_6552 <= 1'h0;
      p14_bit_slice_6553 <= 1'h0;
      p14_bit_slice_6554 <= 1'h0;
      p14_bit_slice_6555 <= 1'h0;
      p14_negated <= 1'h0;
      p15_b <= 32'h0000_0000;
      p15_uge_6629 <= 1'h0;
      p15_bivisor__1 <= 33'h0_0000_0000;
      p15_uge_6637 <= 1'h0;
      p15_uge_6719 <= 1'h0;
      p15_uge_6801 <= 1'h0;
      p15_uge_6881 <= 1'h0;
      p15_uge_6963 <= 1'h0;
      p15_uge_6969 <= 1'h0;
      p15_uge_7049 <= 1'h0;
      p15_uge_7131 <= 1'h0;
      p15_uge_7211 <= 1'h0;
      p15_uge_7293 <= 1'h0;
      p15_uge_7299 <= 1'h0;
      p15_uge_7379 <= 1'h0;
      p15_uge_7461 <= 1'h0;
      p15_uge_7541 <= 1'h0;
      p15_uge_7623 <= 1'h0;
      p15_uge_7629 <= 1'h0;
      p15_uge_7709 <= 1'h0;
      p15_uge_7791 <= 1'h0;
      p15_r__83 <= 32'h0000_0000;
      p15_bit_slice_6543 <= 1'h0;
      p15_bit_slice_6544 <= 1'h0;
      p15_bit_slice_6545 <= 1'h0;
      p15_bit_slice_6546 <= 1'h0;
      p15_bit_slice_6547 <= 1'h0;
      p15_bit_slice_6548 <= 1'h0;
      p15_bit_slice_6549 <= 1'h0;
      p15_bit_slice_6550 <= 1'h0;
      p15_bit_slice_6551 <= 1'h0;
      p15_bit_slice_6552 <= 1'h0;
      p15_bit_slice_6553 <= 1'h0;
      p15_bit_slice_6554 <= 1'h0;
      p15_bit_slice_6555 <= 1'h0;
      p15_negated <= 1'h0;
      p16_b <= 32'h0000_0000;
      p16_uge_6629 <= 1'h0;
      p16_bivisor__1 <= 33'h0_0000_0000;
      p16_uge_6637 <= 1'h0;
      p16_uge_6719 <= 1'h0;
      p16_uge_6801 <= 1'h0;
      p16_uge_6881 <= 1'h0;
      p16_uge_6963 <= 1'h0;
      p16_uge_6969 <= 1'h0;
      p16_uge_7049 <= 1'h0;
      p16_uge_7131 <= 1'h0;
      p16_uge_7211 <= 1'h0;
      p16_uge_7293 <= 1'h0;
      p16_uge_7299 <= 1'h0;
      p16_uge_7379 <= 1'h0;
      p16_uge_7461 <= 1'h0;
      p16_uge_7541 <= 1'h0;
      p16_uge_7623 <= 1'h0;
      p16_uge_7629 <= 1'h0;
      p16_uge_7709 <= 1'h0;
      p16_uge_7791 <= 1'h0;
      p16_uge_7871 <= 1'h0;
      p16_r__84 <= 32'h0000_0000;
      p16_bit_slice_6544 <= 1'h0;
      p16_bit_slice_7874 <= 31'h0000_0000;
      p16_bit_slice_6545 <= 1'h0;
      p16_bit_slice_6546 <= 1'h0;
      p16_bit_slice_6547 <= 1'h0;
      p16_bit_slice_6548 <= 1'h0;
      p16_bit_slice_6549 <= 1'h0;
      p16_bit_slice_6550 <= 1'h0;
      p16_bit_slice_6551 <= 1'h0;
      p16_bit_slice_6552 <= 1'h0;
      p16_bit_slice_6553 <= 1'h0;
      p16_bit_slice_6554 <= 1'h0;
      p16_bit_slice_6555 <= 1'h0;
      p16_negated <= 1'h0;
      p17_b <= 32'h0000_0000;
      p17_uge_6629 <= 1'h0;
      p17_bivisor__1 <= 33'h0_0000_0000;
      p17_uge_6637 <= 1'h0;
      p17_uge_6719 <= 1'h0;
      p17_uge_6801 <= 1'h0;
      p17_uge_6881 <= 1'h0;
      p17_uge_6963 <= 1'h0;
      p17_uge_6969 <= 1'h0;
      p17_uge_7049 <= 1'h0;
      p17_uge_7131 <= 1'h0;
      p17_uge_7211 <= 1'h0;
      p17_uge_7293 <= 1'h0;
      p17_uge_7299 <= 1'h0;
      p17_uge_7379 <= 1'h0;
      p17_uge_7461 <= 1'h0;
      p17_uge_7541 <= 1'h0;
      p17_uge_7623 <= 1'h0;
      p17_uge_7629 <= 1'h0;
      p17_uge_7709 <= 1'h0;
      p17_uge_7791 <= 1'h0;
      p17_uge_7871 <= 1'h0;
      p17_uge_7953 <= 1'h0;
      p17_concat_7958 <= 32'h0000_0000;
      p17_uge_7959 <= 1'h0;
      p17_bit_slice_6546 <= 1'h0;
      p17_bit_slice_6547 <= 1'h0;
      p17_bit_slice_6548 <= 1'h0;
      p17_bit_slice_6549 <= 1'h0;
      p17_bit_slice_6550 <= 1'h0;
      p17_bit_slice_6551 <= 1'h0;
      p17_bit_slice_6552 <= 1'h0;
      p17_bit_slice_6553 <= 1'h0;
      p17_bit_slice_6554 <= 1'h0;
      p17_bit_slice_6555 <= 1'h0;
      p17_negated <= 1'h0;
      p18_b <= 32'h0000_0000;
      p18_uge_6629 <= 1'h0;
      p18_bivisor__1 <= 33'h0_0000_0000;
      p18_uge_6637 <= 1'h0;
      p18_uge_6719 <= 1'h0;
      p18_uge_6801 <= 1'h0;
      p18_uge_6881 <= 1'h0;
      p18_uge_6963 <= 1'h0;
      p18_uge_6969 <= 1'h0;
      p18_uge_7049 <= 1'h0;
      p18_uge_7131 <= 1'h0;
      p18_uge_7211 <= 1'h0;
      p18_uge_7293 <= 1'h0;
      p18_uge_7299 <= 1'h0;
      p18_uge_7379 <= 1'h0;
      p18_uge_7461 <= 1'h0;
      p18_uge_7541 <= 1'h0;
      p18_uge_7623 <= 1'h0;
      p18_uge_7629 <= 1'h0;
      p18_uge_7709 <= 1'h0;
      p18_uge_7791 <= 1'h0;
      p18_uge_7871 <= 1'h0;
      p18_uge_7953 <= 1'h0;
      p18_uge_7959 <= 1'h0;
      p18_concat_8038 <= 32'h0000_0000;
      p18_uge_8039 <= 1'h0;
      p18_sub_8040 <= 32'h0000_0000;
      p18_bit_slice_6547 <= 1'h0;
      p18_bit_slice_6548 <= 1'h0;
      p18_bit_slice_6549 <= 1'h0;
      p18_bit_slice_6550 <= 1'h0;
      p18_bit_slice_6551 <= 1'h0;
      p18_bit_slice_6552 <= 1'h0;
      p18_bit_slice_6553 <= 1'h0;
      p18_bit_slice_6554 <= 1'h0;
      p18_bit_slice_6555 <= 1'h0;
      p18_negated <= 1'h0;
      p19_b <= 32'h0000_0000;
      p19_uge_6629 <= 1'h0;
      p19_bivisor__1 <= 33'h0_0000_0000;
      p19_uge_6637 <= 1'h0;
      p19_uge_6719 <= 1'h0;
      p19_uge_6801 <= 1'h0;
      p19_uge_6881 <= 1'h0;
      p19_uge_6963 <= 1'h0;
      p19_uge_6969 <= 1'h0;
      p19_uge_7049 <= 1'h0;
      p19_uge_7131 <= 1'h0;
      p19_uge_7211 <= 1'h0;
      p19_uge_7293 <= 1'h0;
      p19_uge_7299 <= 1'h0;
      p19_uge_7379 <= 1'h0;
      p19_uge_7461 <= 1'h0;
      p19_uge_7541 <= 1'h0;
      p19_uge_7623 <= 1'h0;
      p19_uge_7629 <= 1'h0;
      p19_uge_7709 <= 1'h0;
      p19_uge_7791 <= 1'h0;
      p19_uge_7871 <= 1'h0;
      p19_uge_7953 <= 1'h0;
      p19_uge_7959 <= 1'h0;
      p19_uge_8039 <= 1'h0;
      p19_uge_8121 <= 1'h0;
      p19_r__88 <= 32'h0000_0000;
      p19_bit_slice_6548 <= 1'h0;
      p19_bit_slice_6549 <= 1'h0;
      p19_bit_slice_6550 <= 1'h0;
      p19_bit_slice_6551 <= 1'h0;
      p19_bit_slice_6552 <= 1'h0;
      p19_bit_slice_6553 <= 1'h0;
      p19_bit_slice_6554 <= 1'h0;
      p19_bit_slice_6555 <= 1'h0;
      p19_negated <= 1'h0;
      p20_b <= 32'h0000_0000;
      p20_uge_6629 <= 1'h0;
      p20_bivisor__1 <= 33'h0_0000_0000;
      p20_uge_6637 <= 1'h0;
      p20_uge_6719 <= 1'h0;
      p20_uge_6801 <= 1'h0;
      p20_uge_6881 <= 1'h0;
      p20_uge_6963 <= 1'h0;
      p20_uge_6969 <= 1'h0;
      p20_uge_7049 <= 1'h0;
      p20_uge_7131 <= 1'h0;
      p20_uge_7211 <= 1'h0;
      p20_uge_7293 <= 1'h0;
      p20_uge_7299 <= 1'h0;
      p20_uge_7379 <= 1'h0;
      p20_uge_7461 <= 1'h0;
      p20_uge_7541 <= 1'h0;
      p20_uge_7623 <= 1'h0;
      p20_uge_7629 <= 1'h0;
      p20_uge_7709 <= 1'h0;
      p20_uge_7791 <= 1'h0;
      p20_uge_7871 <= 1'h0;
      p20_uge_7953 <= 1'h0;
      p20_uge_7959 <= 1'h0;
      p20_uge_8039 <= 1'h0;
      p20_uge_8121 <= 1'h0;
      p20_uge_8201 <= 1'h0;
      p20_r__89 <= 32'h0000_0000;
      p20_bit_slice_6549 <= 1'h0;
      p20_bit_slice_8204 <= 31'h0000_0000;
      p20_bit_slice_6550 <= 1'h0;
      p20_bit_slice_6551 <= 1'h0;
      p20_bit_slice_6552 <= 1'h0;
      p20_bit_slice_6553 <= 1'h0;
      p20_bit_slice_6554 <= 1'h0;
      p20_bit_slice_6555 <= 1'h0;
      p20_negated <= 1'h0;
      p21_b <= 32'h0000_0000;
      p21_uge_6629 <= 1'h0;
      p21_bivisor__1 <= 33'h0_0000_0000;
      p21_uge_6637 <= 1'h0;
      p21_uge_6719 <= 1'h0;
      p21_uge_6801 <= 1'h0;
      p21_uge_6881 <= 1'h0;
      p21_uge_6963 <= 1'h0;
      p21_uge_6969 <= 1'h0;
      p21_uge_7049 <= 1'h0;
      p21_uge_7131 <= 1'h0;
      p21_uge_7211 <= 1'h0;
      p21_uge_7293 <= 1'h0;
      p21_uge_7299 <= 1'h0;
      p21_uge_7379 <= 1'h0;
      p21_uge_7461 <= 1'h0;
      p21_uge_7541 <= 1'h0;
      p21_uge_7623 <= 1'h0;
      p21_uge_7629 <= 1'h0;
      p21_uge_7709 <= 1'h0;
      p21_uge_7791 <= 1'h0;
      p21_uge_7871 <= 1'h0;
      p21_uge_7953 <= 1'h0;
      p21_uge_7959 <= 1'h0;
      p21_uge_8039 <= 1'h0;
      p21_uge_8121 <= 1'h0;
      p21_uge_8201 <= 1'h0;
      p21_uge_8283 <= 1'h0;
      p21_concat_8288 <= 32'h0000_0000;
      p21_uge_8289 <= 1'h0;
      p21_bit_slice_6551 <= 1'h0;
      p21_bit_slice_6552 <= 1'h0;
      p21_bit_slice_6553 <= 1'h0;
      p21_bit_slice_6554 <= 1'h0;
      p21_bit_slice_6555 <= 1'h0;
      p21_negated <= 1'h0;
      p22_b <= 32'h0000_0000;
      p22_uge_6629 <= 1'h0;
      p22_bivisor__1 <= 33'h0_0000_0000;
      p22_uge_6637 <= 1'h0;
      p22_uge_6719 <= 1'h0;
      p22_uge_6801 <= 1'h0;
      p22_uge_6881 <= 1'h0;
      p22_uge_6963 <= 1'h0;
      p22_uge_6969 <= 1'h0;
      p22_uge_7049 <= 1'h0;
      p22_uge_7131 <= 1'h0;
      p22_uge_7211 <= 1'h0;
      p22_uge_7293 <= 1'h0;
      p22_uge_7299 <= 1'h0;
      p22_uge_7379 <= 1'h0;
      p22_uge_7461 <= 1'h0;
      p22_uge_7541 <= 1'h0;
      p22_uge_7623 <= 1'h0;
      p22_uge_7629 <= 1'h0;
      p22_uge_7709 <= 1'h0;
      p22_uge_7791 <= 1'h0;
      p22_uge_7871 <= 1'h0;
      p22_uge_7953 <= 1'h0;
      p22_uge_7959 <= 1'h0;
      p22_uge_8039 <= 1'h0;
      p22_uge_8121 <= 1'h0;
      p22_uge_8201 <= 1'h0;
      p22_uge_8283 <= 1'h0;
      p22_uge_8289 <= 1'h0;
      p22_concat_8368 <= 32'h0000_0000;
      p22_uge_8369 <= 1'h0;
      p22_sub_8370 <= 32'h0000_0000;
      p22_bit_slice_6552 <= 1'h0;
      p22_bit_slice_6553 <= 1'h0;
      p22_bit_slice_6554 <= 1'h0;
      p22_bit_slice_6555 <= 1'h0;
      p22_negated <= 1'h0;
      p23_b <= 32'h0000_0000;
      p23_uge_6629 <= 1'h0;
      p23_bivisor__1 <= 33'h0_0000_0000;
      p23_uge_6637 <= 1'h0;
      p23_uge_6719 <= 1'h0;
      p23_uge_6801 <= 1'h0;
      p23_uge_6881 <= 1'h0;
      p23_uge_6963 <= 1'h0;
      p23_uge_6969 <= 1'h0;
      p23_uge_7049 <= 1'h0;
      p23_uge_7131 <= 1'h0;
      p23_uge_7211 <= 1'h0;
      p23_uge_7293 <= 1'h0;
      p23_uge_7299 <= 1'h0;
      p23_uge_7379 <= 1'h0;
      p23_uge_7461 <= 1'h0;
      p23_uge_7541 <= 1'h0;
      p23_uge_7623 <= 1'h0;
      p23_uge_7629 <= 1'h0;
      p23_uge_7709 <= 1'h0;
      p23_uge_7791 <= 1'h0;
      p23_uge_7871 <= 1'h0;
      p23_uge_7953 <= 1'h0;
      p23_uge_7959 <= 1'h0;
      p23_uge_8039 <= 1'h0;
      p23_uge_8121 <= 1'h0;
      p23_uge_8201 <= 1'h0;
      p23_uge_8283 <= 1'h0;
      p23_uge_8289 <= 1'h0;
      p23_uge_8369 <= 1'h0;
      p23_uge_8451 <= 1'h0;
      p23_r__93 <= 32'h0000_0000;
      p23_bit_slice_6553 <= 1'h0;
      p23_bit_slice_6554 <= 1'h0;
      p23_bit_slice_6555 <= 1'h0;
      p23_negated <= 1'h0;
      p24_b <= 32'h0000_0000;
      p24_uge_6629 <= 1'h0;
      p24_bivisor__1 <= 33'h0_0000_0000;
      p24_uge_6637 <= 1'h0;
      p24_uge_6719 <= 1'h0;
      p24_uge_6801 <= 1'h0;
      p24_uge_6881 <= 1'h0;
      p24_uge_6963 <= 1'h0;
      p24_uge_6969 <= 1'h0;
      p24_uge_7049 <= 1'h0;
      p24_uge_7131 <= 1'h0;
      p24_uge_7211 <= 1'h0;
      p24_uge_7293 <= 1'h0;
      p24_uge_7299 <= 1'h0;
      p24_uge_7379 <= 1'h0;
      p24_uge_7461 <= 1'h0;
      p24_uge_7541 <= 1'h0;
      p24_uge_7623 <= 1'h0;
      p24_uge_7629 <= 1'h0;
      p24_uge_7709 <= 1'h0;
      p24_uge_7791 <= 1'h0;
      p24_uge_7871 <= 1'h0;
      p24_uge_7953 <= 1'h0;
      p24_uge_7959 <= 1'h0;
      p24_uge_8039 <= 1'h0;
      p24_uge_8121 <= 1'h0;
      p24_uge_8201 <= 1'h0;
      p24_uge_8283 <= 1'h0;
      p24_uge_8289 <= 1'h0;
      p24_uge_8369 <= 1'h0;
      p24_uge_8451 <= 1'h0;
      p24_uge_8531 <= 1'h0;
      p24_r__94 <= 32'h0000_0000;
      p24_bit_slice_6554 <= 1'h0;
      p24_bit_slice_8534 <= 31'h0000_0000;
      p24_bit_slice_6555 <= 1'h0;
      p24_negated <= 1'h0;
      p25_uge_6629 <= 1'h0;
      p25_uge_6637 <= 1'h0;
      p25_uge_6719 <= 1'h0;
      p25_uge_6801 <= 1'h0;
      p25_uge_6881 <= 1'h0;
      p25_uge_6963 <= 1'h0;
      p25_uge_6969 <= 1'h0;
      p25_uge_7049 <= 1'h0;
      p25_uge_7131 <= 1'h0;
      p25_uge_7211 <= 1'h0;
      p25_uge_7293 <= 1'h0;
      p25_uge_7299 <= 1'h0;
      p25_uge_7379 <= 1'h0;
      p25_uge_7461 <= 1'h0;
      p25_uge_7541 <= 1'h0;
      p25_uge_7623 <= 1'h0;
      p25_uge_7629 <= 1'h0;
      p25_uge_7709 <= 1'h0;
      p25_uge_7791 <= 1'h0;
      p25_uge_7871 <= 1'h0;
      p25_uge_7953 <= 1'h0;
      p25_uge_7959 <= 1'h0;
      p25_uge_8039 <= 1'h0;
      p25_uge_8121 <= 1'h0;
      p25_uge_8201 <= 1'h0;
      p25_uge_8283 <= 1'h0;
      p25_uge_8289 <= 1'h0;
      p25_uge_8369 <= 1'h0;
      p25_uge_8451 <= 1'h0;
      p25_uge_8531 <= 1'h0;
      p25_uge_8613 <= 1'h0;
      p25_q__32_squeezed_portion_0_width_1 <= 1'h0;
      p25_negated <= 1'h0;
      p0_valid <= 1'h0;
      p1_valid <= 1'h0;
      p2_valid <= 1'h0;
      p3_valid <= 1'h0;
      p4_valid <= 1'h0;
      p5_valid <= 1'h0;
      p6_valid <= 1'h0;
      p7_valid <= 1'h0;
      p8_valid <= 1'h0;
      p9_valid <= 1'h0;
      p10_valid <= 1'h0;
      p11_valid <= 1'h0;
      p12_valid <= 1'h0;
      p13_valid <= 1'h0;
      p14_valid <= 1'h0;
      p15_valid <= 1'h0;
      p16_valid <= 1'h0;
      p17_valid <= 1'h0;
      p18_valid <= 1'h0;
      p19_valid <= 1'h0;
      p20_valid <= 1'h0;
      p21_valid <= 1'h0;
      p22_valid <= 1'h0;
      p23_valid <= 1'h0;
      p24_valid <= 1'h0;
      p25_valid <= 1'h0;
      p26_valid <= 1'h0;
      p27_valid <= 1'h0;
      p28_valid <= 1'h0;
      p29_valid <= 1'h0;
      p30_valid <= 1'h0;
      lhs_reg <= 32'h0000_0000;
      lhs_valid_reg <= 1'h0;
      rhs_reg <= 32'h0000_0000;
      rhs_valid_reg <= 1'h0;
      result_reg <= 32'h0000_0000;
      result_valid_reg <= 1'h0;
    end else begin
      p0_sign_a <= p0_data_enable ? sign_a : p0_sign_a;
      p0_b <= p0_data_enable ? rhs_reg : p0_b;
      p0_bit_slice_6525 <= p0_data_enable ? bit_slice_6525 : p0_bit_slice_6525;
      p0_bit_slice_6526 <= p0_data_enable ? bit_slice_6526 : p0_bit_slice_6526;
      p0_bit_slice_6527 <= p0_data_enable ? bit_slice_6527 : p0_bit_slice_6527;
      p0_bit_slice_6528 <= p0_data_enable ? bit_slice_6528 : p0_bit_slice_6528;
      p0_bit_slice_6529 <= p0_data_enable ? bit_slice_6529 : p0_bit_slice_6529;
      p0_bit_slice_6530 <= p0_data_enable ? bit_slice_6530 : p0_bit_slice_6530;
      p0_bit_slice_6531 <= p0_data_enable ? bit_slice_6531 : p0_bit_slice_6531;
      p0_bit_slice_6532 <= p0_data_enable ? bit_slice_6532 : p0_bit_slice_6532;
      p0_bit_slice_6533 <= p0_data_enable ? bit_slice_6533 : p0_bit_slice_6533;
      p0_bit_slice_6534 <= p0_data_enable ? bit_slice_6534 : p0_bit_slice_6534;
      p0_bit_slice_6535 <= p0_data_enable ? bit_slice_6535 : p0_bit_slice_6535;
      p0_bit_slice_6536 <= p0_data_enable ? bit_slice_6536 : p0_bit_slice_6536;
      p0_bit_slice_6537 <= p0_data_enable ? bit_slice_6537 : p0_bit_slice_6537;
      p0_bit_slice_6538 <= p0_data_enable ? bit_slice_6538 : p0_bit_slice_6538;
      p0_bit_slice_6539 <= p0_data_enable ? bit_slice_6539 : p0_bit_slice_6539;
      p0_bit_slice_6540 <= p0_data_enable ? bit_slice_6540 : p0_bit_slice_6540;
      p0_bit_slice_6541 <= p0_data_enable ? bit_slice_6541 : p0_bit_slice_6541;
      p0_bit_slice_6542 <= p0_data_enable ? bit_slice_6542 : p0_bit_slice_6542;
      p0_bit_slice_6543 <= p0_data_enable ? bit_slice_6543 : p0_bit_slice_6543;
      p0_bit_slice_6544 <= p0_data_enable ? bit_slice_6544 : p0_bit_slice_6544;
      p0_bit_slice_6545 <= p0_data_enable ? bit_slice_6545 : p0_bit_slice_6545;
      p0_bit_slice_6546 <= p0_data_enable ? bit_slice_6546 : p0_bit_slice_6546;
      p0_bit_slice_6547 <= p0_data_enable ? bit_slice_6547 : p0_bit_slice_6547;
      p0_bit_slice_6548 <= p0_data_enable ? bit_slice_6548 : p0_bit_slice_6548;
      p0_bit_slice_6549 <= p0_data_enable ? bit_slice_6549 : p0_bit_slice_6549;
      p0_bit_slice_6550 <= p0_data_enable ? bit_slice_6550 : p0_bit_slice_6550;
      p0_bit_slice_6551 <= p0_data_enable ? bit_slice_6551 : p0_bit_slice_6551;
      p0_bit_slice_6552 <= p0_data_enable ? bit_slice_6552 : p0_bit_slice_6552;
      p0_bit_slice_6553 <= p0_data_enable ? bit_slice_6553 : p0_bit_slice_6553;
      p0_bit_slice_6554 <= p0_data_enable ? bit_slice_6554 : p0_bit_slice_6554;
      p0_bit_slice_6555 <= p0_data_enable ? bit_slice_6555 : p0_bit_slice_6555;
      p1_b <= p1_data_enable ? p0_b : p1_b;
      p1_uge_6629 <= p1_data_enable ? uge_6629 : p1_uge_6629;
      p1_bivisor__1 <= p1_data_enable ? bivisor__1 : p1_bivisor__1;
      p1_concat_6636 <= p1_data_enable ? concat_6636 : p1_concat_6636;
      p1_uge_6637 <= p1_data_enable ? uge_6637 : p1_uge_6637;
      p1_bit_slice_6526 <= p1_data_enable ? p0_bit_slice_6526 : p1_bit_slice_6526;
      p1_bit_slice_6527 <= p1_data_enable ? p0_bit_slice_6527 : p1_bit_slice_6527;
      p1_bit_slice_6528 <= p1_data_enable ? p0_bit_slice_6528 : p1_bit_slice_6528;
      p1_bit_slice_6529 <= p1_data_enable ? p0_bit_slice_6529 : p1_bit_slice_6529;
      p1_bit_slice_6530 <= p1_data_enable ? p0_bit_slice_6530 : p1_bit_slice_6530;
      p1_bit_slice_6531 <= p1_data_enable ? p0_bit_slice_6531 : p1_bit_slice_6531;
      p1_bit_slice_6532 <= p1_data_enable ? p0_bit_slice_6532 : p1_bit_slice_6532;
      p1_bit_slice_6533 <= p1_data_enable ? p0_bit_slice_6533 : p1_bit_slice_6533;
      p1_bit_slice_6534 <= p1_data_enable ? p0_bit_slice_6534 : p1_bit_slice_6534;
      p1_bit_slice_6535 <= p1_data_enable ? p0_bit_slice_6535 : p1_bit_slice_6535;
      p1_bit_slice_6536 <= p1_data_enable ? p0_bit_slice_6536 : p1_bit_slice_6536;
      p1_bit_slice_6537 <= p1_data_enable ? p0_bit_slice_6537 : p1_bit_slice_6537;
      p1_bit_slice_6538 <= p1_data_enable ? p0_bit_slice_6538 : p1_bit_slice_6538;
      p1_bit_slice_6539 <= p1_data_enable ? p0_bit_slice_6539 : p1_bit_slice_6539;
      p1_bit_slice_6540 <= p1_data_enable ? p0_bit_slice_6540 : p1_bit_slice_6540;
      p1_bit_slice_6541 <= p1_data_enable ? p0_bit_slice_6541 : p1_bit_slice_6541;
      p1_bit_slice_6542 <= p1_data_enable ? p0_bit_slice_6542 : p1_bit_slice_6542;
      p1_bit_slice_6543 <= p1_data_enable ? p0_bit_slice_6543 : p1_bit_slice_6543;
      p1_bit_slice_6544 <= p1_data_enable ? p0_bit_slice_6544 : p1_bit_slice_6544;
      p1_bit_slice_6545 <= p1_data_enable ? p0_bit_slice_6545 : p1_bit_slice_6545;
      p1_bit_slice_6546 <= p1_data_enable ? p0_bit_slice_6546 : p1_bit_slice_6546;
      p1_bit_slice_6547 <= p1_data_enable ? p0_bit_slice_6547 : p1_bit_slice_6547;
      p1_bit_slice_6548 <= p1_data_enable ? p0_bit_slice_6548 : p1_bit_slice_6548;
      p1_bit_slice_6549 <= p1_data_enable ? p0_bit_slice_6549 : p1_bit_slice_6549;
      p1_bit_slice_6550 <= p1_data_enable ? p0_bit_slice_6550 : p1_bit_slice_6550;
      p1_bit_slice_6551 <= p1_data_enable ? p0_bit_slice_6551 : p1_bit_slice_6551;
      p1_bit_slice_6552 <= p1_data_enable ? p0_bit_slice_6552 : p1_bit_slice_6552;
      p1_bit_slice_6553 <= p1_data_enable ? p0_bit_slice_6553 : p1_bit_slice_6553;
      p1_bit_slice_6554 <= p1_data_enable ? p0_bit_slice_6554 : p1_bit_slice_6554;
      p1_bit_slice_6555 <= p1_data_enable ? p0_bit_slice_6555 : p1_bit_slice_6555;
      p1_negated <= p1_data_enable ? negated : p1_negated;
      p2_b <= p2_data_enable ? p1_b : p2_b;
      p2_uge_6629 <= p2_data_enable ? p1_uge_6629 : p2_uge_6629;
      p2_bivisor__1 <= p2_data_enable ? p1_bivisor__1 : p2_bivisor__1;
      p2_uge_6637 <= p2_data_enable ? p1_uge_6637 : p2_uge_6637;
      p2_concat_6718 <= p2_data_enable ? concat_6718 : p2_concat_6718;
      p2_uge_6719 <= p2_data_enable ? uge_6719 : p2_uge_6719;
      p2_sub_6720 <= p2_data_enable ? sub_6720 : p2_sub_6720;
      p2_bit_slice_6527 <= p2_data_enable ? p1_bit_slice_6527 : p2_bit_slice_6527;
      p2_bit_slice_6528 <= p2_data_enable ? p1_bit_slice_6528 : p2_bit_slice_6528;
      p2_bit_slice_6529 <= p2_data_enable ? p1_bit_slice_6529 : p2_bit_slice_6529;
      p2_bit_slice_6530 <= p2_data_enable ? p1_bit_slice_6530 : p2_bit_slice_6530;
      p2_bit_slice_6531 <= p2_data_enable ? p1_bit_slice_6531 : p2_bit_slice_6531;
      p2_bit_slice_6532 <= p2_data_enable ? p1_bit_slice_6532 : p2_bit_slice_6532;
      p2_bit_slice_6533 <= p2_data_enable ? p1_bit_slice_6533 : p2_bit_slice_6533;
      p2_bit_slice_6534 <= p2_data_enable ? p1_bit_slice_6534 : p2_bit_slice_6534;
      p2_bit_slice_6535 <= p2_data_enable ? p1_bit_slice_6535 : p2_bit_slice_6535;
      p2_bit_slice_6536 <= p2_data_enable ? p1_bit_slice_6536 : p2_bit_slice_6536;
      p2_bit_slice_6537 <= p2_data_enable ? p1_bit_slice_6537 : p2_bit_slice_6537;
      p2_bit_slice_6538 <= p2_data_enable ? p1_bit_slice_6538 : p2_bit_slice_6538;
      p2_bit_slice_6539 <= p2_data_enable ? p1_bit_slice_6539 : p2_bit_slice_6539;
      p2_bit_slice_6540 <= p2_data_enable ? p1_bit_slice_6540 : p2_bit_slice_6540;
      p2_bit_slice_6541 <= p2_data_enable ? p1_bit_slice_6541 : p2_bit_slice_6541;
      p2_bit_slice_6542 <= p2_data_enable ? p1_bit_slice_6542 : p2_bit_slice_6542;
      p2_bit_slice_6543 <= p2_data_enable ? p1_bit_slice_6543 : p2_bit_slice_6543;
      p2_bit_slice_6544 <= p2_data_enable ? p1_bit_slice_6544 : p2_bit_slice_6544;
      p2_bit_slice_6545 <= p2_data_enable ? p1_bit_slice_6545 : p2_bit_slice_6545;
      p2_bit_slice_6546 <= p2_data_enable ? p1_bit_slice_6546 : p2_bit_slice_6546;
      p2_bit_slice_6547 <= p2_data_enable ? p1_bit_slice_6547 : p2_bit_slice_6547;
      p2_bit_slice_6548 <= p2_data_enable ? p1_bit_slice_6548 : p2_bit_slice_6548;
      p2_bit_slice_6549 <= p2_data_enable ? p1_bit_slice_6549 : p2_bit_slice_6549;
      p2_bit_slice_6550 <= p2_data_enable ? p1_bit_slice_6550 : p2_bit_slice_6550;
      p2_bit_slice_6551 <= p2_data_enable ? p1_bit_slice_6551 : p2_bit_slice_6551;
      p2_bit_slice_6552 <= p2_data_enable ? p1_bit_slice_6552 : p2_bit_slice_6552;
      p2_bit_slice_6553 <= p2_data_enable ? p1_bit_slice_6553 : p2_bit_slice_6553;
      p2_bit_slice_6554 <= p2_data_enable ? p1_bit_slice_6554 : p2_bit_slice_6554;
      p2_bit_slice_6555 <= p2_data_enable ? p1_bit_slice_6555 : p2_bit_slice_6555;
      p2_negated <= p2_data_enable ? p1_negated : p2_negated;
      p3_b <= p3_data_enable ? p2_b : p3_b;
      p3_uge_6629 <= p3_data_enable ? p2_uge_6629 : p3_uge_6629;
      p3_bivisor__1 <= p3_data_enable ? p2_bivisor__1 : p3_bivisor__1;
      p3_uge_6637 <= p3_data_enable ? p2_uge_6637 : p3_uge_6637;
      p3_uge_6719 <= p3_data_enable ? p2_uge_6719 : p3_uge_6719;
      p3_uge_6801 <= p3_data_enable ? uge_6801 : p3_uge_6801;
      p3_r__68 <= p3_data_enable ? r__68 : p3_r__68;
      p3_bit_slice_6528 <= p3_data_enable ? p2_bit_slice_6528 : p3_bit_slice_6528;
      p3_bit_slice_6529 <= p3_data_enable ? p2_bit_slice_6529 : p3_bit_slice_6529;
      p3_bit_slice_6530 <= p3_data_enable ? p2_bit_slice_6530 : p3_bit_slice_6530;
      p3_bit_slice_6531 <= p3_data_enable ? p2_bit_slice_6531 : p3_bit_slice_6531;
      p3_bit_slice_6532 <= p3_data_enable ? p2_bit_slice_6532 : p3_bit_slice_6532;
      p3_bit_slice_6533 <= p3_data_enable ? p2_bit_slice_6533 : p3_bit_slice_6533;
      p3_bit_slice_6534 <= p3_data_enable ? p2_bit_slice_6534 : p3_bit_slice_6534;
      p3_bit_slice_6535 <= p3_data_enable ? p2_bit_slice_6535 : p3_bit_slice_6535;
      p3_bit_slice_6536 <= p3_data_enable ? p2_bit_slice_6536 : p3_bit_slice_6536;
      p3_bit_slice_6537 <= p3_data_enable ? p2_bit_slice_6537 : p3_bit_slice_6537;
      p3_bit_slice_6538 <= p3_data_enable ? p2_bit_slice_6538 : p3_bit_slice_6538;
      p3_bit_slice_6539 <= p3_data_enable ? p2_bit_slice_6539 : p3_bit_slice_6539;
      p3_bit_slice_6540 <= p3_data_enable ? p2_bit_slice_6540 : p3_bit_slice_6540;
      p3_bit_slice_6541 <= p3_data_enable ? p2_bit_slice_6541 : p3_bit_slice_6541;
      p3_bit_slice_6542 <= p3_data_enable ? p2_bit_slice_6542 : p3_bit_slice_6542;
      p3_bit_slice_6543 <= p3_data_enable ? p2_bit_slice_6543 : p3_bit_slice_6543;
      p3_bit_slice_6544 <= p3_data_enable ? p2_bit_slice_6544 : p3_bit_slice_6544;
      p3_bit_slice_6545 <= p3_data_enable ? p2_bit_slice_6545 : p3_bit_slice_6545;
      p3_bit_slice_6546 <= p3_data_enable ? p2_bit_slice_6546 : p3_bit_slice_6546;
      p3_bit_slice_6547 <= p3_data_enable ? p2_bit_slice_6547 : p3_bit_slice_6547;
      p3_bit_slice_6548 <= p3_data_enable ? p2_bit_slice_6548 : p3_bit_slice_6548;
      p3_bit_slice_6549 <= p3_data_enable ? p2_bit_slice_6549 : p3_bit_slice_6549;
      p3_bit_slice_6550 <= p3_data_enable ? p2_bit_slice_6550 : p3_bit_slice_6550;
      p3_bit_slice_6551 <= p3_data_enable ? p2_bit_slice_6551 : p3_bit_slice_6551;
      p3_bit_slice_6552 <= p3_data_enable ? p2_bit_slice_6552 : p3_bit_slice_6552;
      p3_bit_slice_6553 <= p3_data_enable ? p2_bit_slice_6553 : p3_bit_slice_6553;
      p3_bit_slice_6554 <= p3_data_enable ? p2_bit_slice_6554 : p3_bit_slice_6554;
      p3_bit_slice_6555 <= p3_data_enable ? p2_bit_slice_6555 : p3_bit_slice_6555;
      p3_negated <= p3_data_enable ? p2_negated : p3_negated;
      p4_b <= p4_data_enable ? p3_b : p4_b;
      p4_uge_6629 <= p4_data_enable ? p3_uge_6629 : p4_uge_6629;
      p4_bivisor__1 <= p4_data_enable ? p3_bivisor__1 : p4_bivisor__1;
      p4_uge_6637 <= p4_data_enable ? p3_uge_6637 : p4_uge_6637;
      p4_uge_6719 <= p4_data_enable ? p3_uge_6719 : p4_uge_6719;
      p4_uge_6801 <= p4_data_enable ? p3_uge_6801 : p4_uge_6801;
      p4_uge_6881 <= p4_data_enable ? uge_6881 : p4_uge_6881;
      p4_r__69 <= p4_data_enable ? r__69 : p4_r__69;
      p4_bit_slice_6529 <= p4_data_enable ? p3_bit_slice_6529 : p4_bit_slice_6529;
      p4_bit_slice_6884 <= p4_data_enable ? bit_slice_6884 : p4_bit_slice_6884;
      p4_bit_slice_6530 <= p4_data_enable ? p3_bit_slice_6530 : p4_bit_slice_6530;
      p4_bit_slice_6531 <= p4_data_enable ? p3_bit_slice_6531 : p4_bit_slice_6531;
      p4_bit_slice_6532 <= p4_data_enable ? p3_bit_slice_6532 : p4_bit_slice_6532;
      p4_bit_slice_6533 <= p4_data_enable ? p3_bit_slice_6533 : p4_bit_slice_6533;
      p4_bit_slice_6534 <= p4_data_enable ? p3_bit_slice_6534 : p4_bit_slice_6534;
      p4_bit_slice_6535 <= p4_data_enable ? p3_bit_slice_6535 : p4_bit_slice_6535;
      p4_bit_slice_6536 <= p4_data_enable ? p3_bit_slice_6536 : p4_bit_slice_6536;
      p4_bit_slice_6537 <= p4_data_enable ? p3_bit_slice_6537 : p4_bit_slice_6537;
      p4_bit_slice_6538 <= p4_data_enable ? p3_bit_slice_6538 : p4_bit_slice_6538;
      p4_bit_slice_6539 <= p4_data_enable ? p3_bit_slice_6539 : p4_bit_slice_6539;
      p4_bit_slice_6540 <= p4_data_enable ? p3_bit_slice_6540 : p4_bit_slice_6540;
      p4_bit_slice_6541 <= p4_data_enable ? p3_bit_slice_6541 : p4_bit_slice_6541;
      p4_bit_slice_6542 <= p4_data_enable ? p3_bit_slice_6542 : p4_bit_slice_6542;
      p4_bit_slice_6543 <= p4_data_enable ? p3_bit_slice_6543 : p4_bit_slice_6543;
      p4_bit_slice_6544 <= p4_data_enable ? p3_bit_slice_6544 : p4_bit_slice_6544;
      p4_bit_slice_6545 <= p4_data_enable ? p3_bit_slice_6545 : p4_bit_slice_6545;
      p4_bit_slice_6546 <= p4_data_enable ? p3_bit_slice_6546 : p4_bit_slice_6546;
      p4_bit_slice_6547 <= p4_data_enable ? p3_bit_slice_6547 : p4_bit_slice_6547;
      p4_bit_slice_6548 <= p4_data_enable ? p3_bit_slice_6548 : p4_bit_slice_6548;
      p4_bit_slice_6549 <= p4_data_enable ? p3_bit_slice_6549 : p4_bit_slice_6549;
      p4_bit_slice_6550 <= p4_data_enable ? p3_bit_slice_6550 : p4_bit_slice_6550;
      p4_bit_slice_6551 <= p4_data_enable ? p3_bit_slice_6551 : p4_bit_slice_6551;
      p4_bit_slice_6552 <= p4_data_enable ? p3_bit_slice_6552 : p4_bit_slice_6552;
      p4_bit_slice_6553 <= p4_data_enable ? p3_bit_slice_6553 : p4_bit_slice_6553;
      p4_bit_slice_6554 <= p4_data_enable ? p3_bit_slice_6554 : p4_bit_slice_6554;
      p4_bit_slice_6555 <= p4_data_enable ? p3_bit_slice_6555 : p4_bit_slice_6555;
      p4_negated <= p4_data_enable ? p3_negated : p4_negated;
      p5_b <= p5_data_enable ? p4_b : p5_b;
      p5_uge_6629 <= p5_data_enable ? p4_uge_6629 : p5_uge_6629;
      p5_bivisor__1 <= p5_data_enable ? p4_bivisor__1 : p5_bivisor__1;
      p5_uge_6637 <= p5_data_enable ? p4_uge_6637 : p5_uge_6637;
      p5_uge_6719 <= p5_data_enable ? p4_uge_6719 : p5_uge_6719;
      p5_uge_6801 <= p5_data_enable ? p4_uge_6801 : p5_uge_6801;
      p5_uge_6881 <= p5_data_enable ? p4_uge_6881 : p5_uge_6881;
      p5_uge_6963 <= p5_data_enable ? uge_6963 : p5_uge_6963;
      p5_concat_6968 <= p5_data_enable ? concat_6968 : p5_concat_6968;
      p5_uge_6969 <= p5_data_enable ? uge_6969 : p5_uge_6969;
      p5_bit_slice_6531 <= p5_data_enable ? p4_bit_slice_6531 : p5_bit_slice_6531;
      p5_bit_slice_6532 <= p5_data_enable ? p4_bit_slice_6532 : p5_bit_slice_6532;
      p5_bit_slice_6533 <= p5_data_enable ? p4_bit_slice_6533 : p5_bit_slice_6533;
      p5_bit_slice_6534 <= p5_data_enable ? p4_bit_slice_6534 : p5_bit_slice_6534;
      p5_bit_slice_6535 <= p5_data_enable ? p4_bit_slice_6535 : p5_bit_slice_6535;
      p5_bit_slice_6536 <= p5_data_enable ? p4_bit_slice_6536 : p5_bit_slice_6536;
      p5_bit_slice_6537 <= p5_data_enable ? p4_bit_slice_6537 : p5_bit_slice_6537;
      p5_bit_slice_6538 <= p5_data_enable ? p4_bit_slice_6538 : p5_bit_slice_6538;
      p5_bit_slice_6539 <= p5_data_enable ? p4_bit_slice_6539 : p5_bit_slice_6539;
      p5_bit_slice_6540 <= p5_data_enable ? p4_bit_slice_6540 : p5_bit_slice_6540;
      p5_bit_slice_6541 <= p5_data_enable ? p4_bit_slice_6541 : p5_bit_slice_6541;
      p5_bit_slice_6542 <= p5_data_enable ? p4_bit_slice_6542 : p5_bit_slice_6542;
      p5_bit_slice_6543 <= p5_data_enable ? p4_bit_slice_6543 : p5_bit_slice_6543;
      p5_bit_slice_6544 <= p5_data_enable ? p4_bit_slice_6544 : p5_bit_slice_6544;
      p5_bit_slice_6545 <= p5_data_enable ? p4_bit_slice_6545 : p5_bit_slice_6545;
      p5_bit_slice_6546 <= p5_data_enable ? p4_bit_slice_6546 : p5_bit_slice_6546;
      p5_bit_slice_6547 <= p5_data_enable ? p4_bit_slice_6547 : p5_bit_slice_6547;
      p5_bit_slice_6548 <= p5_data_enable ? p4_bit_slice_6548 : p5_bit_slice_6548;
      p5_bit_slice_6549 <= p5_data_enable ? p4_bit_slice_6549 : p5_bit_slice_6549;
      p5_bit_slice_6550 <= p5_data_enable ? p4_bit_slice_6550 : p5_bit_slice_6550;
      p5_bit_slice_6551 <= p5_data_enable ? p4_bit_slice_6551 : p5_bit_slice_6551;
      p5_bit_slice_6552 <= p5_data_enable ? p4_bit_slice_6552 : p5_bit_slice_6552;
      p5_bit_slice_6553 <= p5_data_enable ? p4_bit_slice_6553 : p5_bit_slice_6553;
      p5_bit_slice_6554 <= p5_data_enable ? p4_bit_slice_6554 : p5_bit_slice_6554;
      p5_bit_slice_6555 <= p5_data_enable ? p4_bit_slice_6555 : p5_bit_slice_6555;
      p5_negated <= p5_data_enable ? p4_negated : p5_negated;
      p6_b <= p6_data_enable ? p5_b : p6_b;
      p6_uge_6629 <= p6_data_enable ? p5_uge_6629 : p6_uge_6629;
      p6_bivisor__1 <= p6_data_enable ? p5_bivisor__1 : p6_bivisor__1;
      p6_uge_6637 <= p6_data_enable ? p5_uge_6637 : p6_uge_6637;
      p6_uge_6719 <= p6_data_enable ? p5_uge_6719 : p6_uge_6719;
      p6_uge_6801 <= p6_data_enable ? p5_uge_6801 : p6_uge_6801;
      p6_uge_6881 <= p6_data_enable ? p5_uge_6881 : p6_uge_6881;
      p6_uge_6963 <= p6_data_enable ? p5_uge_6963 : p6_uge_6963;
      p6_uge_6969 <= p6_data_enable ? p5_uge_6969 : p6_uge_6969;
      p6_concat_7048 <= p6_data_enable ? concat_7048 : p6_concat_7048;
      p6_uge_7049 <= p6_data_enable ? uge_7049 : p6_uge_7049;
      p6_sub_7050 <= p6_data_enable ? sub_7050 : p6_sub_7050;
      p6_bit_slice_6532 <= p6_data_enable ? p5_bit_slice_6532 : p6_bit_slice_6532;
      p6_bit_slice_6533 <= p6_data_enable ? p5_bit_slice_6533 : p6_bit_slice_6533;
      p6_bit_slice_6534 <= p6_data_enable ? p5_bit_slice_6534 : p6_bit_slice_6534;
      p6_bit_slice_6535 <= p6_data_enable ? p5_bit_slice_6535 : p6_bit_slice_6535;
      p6_bit_slice_6536 <= p6_data_enable ? p5_bit_slice_6536 : p6_bit_slice_6536;
      p6_bit_slice_6537 <= p6_data_enable ? p5_bit_slice_6537 : p6_bit_slice_6537;
      p6_bit_slice_6538 <= p6_data_enable ? p5_bit_slice_6538 : p6_bit_slice_6538;
      p6_bit_slice_6539 <= p6_data_enable ? p5_bit_slice_6539 : p6_bit_slice_6539;
      p6_bit_slice_6540 <= p6_data_enable ? p5_bit_slice_6540 : p6_bit_slice_6540;
      p6_bit_slice_6541 <= p6_data_enable ? p5_bit_slice_6541 : p6_bit_slice_6541;
      p6_bit_slice_6542 <= p6_data_enable ? p5_bit_slice_6542 : p6_bit_slice_6542;
      p6_bit_slice_6543 <= p6_data_enable ? p5_bit_slice_6543 : p6_bit_slice_6543;
      p6_bit_slice_6544 <= p6_data_enable ? p5_bit_slice_6544 : p6_bit_slice_6544;
      p6_bit_slice_6545 <= p6_data_enable ? p5_bit_slice_6545 : p6_bit_slice_6545;
      p6_bit_slice_6546 <= p6_data_enable ? p5_bit_slice_6546 : p6_bit_slice_6546;
      p6_bit_slice_6547 <= p6_data_enable ? p5_bit_slice_6547 : p6_bit_slice_6547;
      p6_bit_slice_6548 <= p6_data_enable ? p5_bit_slice_6548 : p6_bit_slice_6548;
      p6_bit_slice_6549 <= p6_data_enable ? p5_bit_slice_6549 : p6_bit_slice_6549;
      p6_bit_slice_6550 <= p6_data_enable ? p5_bit_slice_6550 : p6_bit_slice_6550;
      p6_bit_slice_6551 <= p6_data_enable ? p5_bit_slice_6551 : p6_bit_slice_6551;
      p6_bit_slice_6552 <= p6_data_enable ? p5_bit_slice_6552 : p6_bit_slice_6552;
      p6_bit_slice_6553 <= p6_data_enable ? p5_bit_slice_6553 : p6_bit_slice_6553;
      p6_bit_slice_6554 <= p6_data_enable ? p5_bit_slice_6554 : p6_bit_slice_6554;
      p6_bit_slice_6555 <= p6_data_enable ? p5_bit_slice_6555 : p6_bit_slice_6555;
      p6_negated <= p6_data_enable ? p5_negated : p6_negated;
      p7_b <= p7_data_enable ? p6_b : p7_b;
      p7_uge_6629 <= p7_data_enable ? p6_uge_6629 : p7_uge_6629;
      p7_bivisor__1 <= p7_data_enable ? p6_bivisor__1 : p7_bivisor__1;
      p7_uge_6637 <= p7_data_enable ? p6_uge_6637 : p7_uge_6637;
      p7_uge_6719 <= p7_data_enable ? p6_uge_6719 : p7_uge_6719;
      p7_uge_6801 <= p7_data_enable ? p6_uge_6801 : p7_uge_6801;
      p7_uge_6881 <= p7_data_enable ? p6_uge_6881 : p7_uge_6881;
      p7_uge_6963 <= p7_data_enable ? p6_uge_6963 : p7_uge_6963;
      p7_uge_6969 <= p7_data_enable ? p6_uge_6969 : p7_uge_6969;
      p7_uge_7049 <= p7_data_enable ? p6_uge_7049 : p7_uge_7049;
      p7_uge_7131 <= p7_data_enable ? uge_7131 : p7_uge_7131;
      p7_r__73 <= p7_data_enable ? r__73 : p7_r__73;
      p7_bit_slice_6533 <= p7_data_enable ? p6_bit_slice_6533 : p7_bit_slice_6533;
      p7_bit_slice_6534 <= p7_data_enable ? p6_bit_slice_6534 : p7_bit_slice_6534;
      p7_bit_slice_6535 <= p7_data_enable ? p6_bit_slice_6535 : p7_bit_slice_6535;
      p7_bit_slice_6536 <= p7_data_enable ? p6_bit_slice_6536 : p7_bit_slice_6536;
      p7_bit_slice_6537 <= p7_data_enable ? p6_bit_slice_6537 : p7_bit_slice_6537;
      p7_bit_slice_6538 <= p7_data_enable ? p6_bit_slice_6538 : p7_bit_slice_6538;
      p7_bit_slice_6539 <= p7_data_enable ? p6_bit_slice_6539 : p7_bit_slice_6539;
      p7_bit_slice_6540 <= p7_data_enable ? p6_bit_slice_6540 : p7_bit_slice_6540;
      p7_bit_slice_6541 <= p7_data_enable ? p6_bit_slice_6541 : p7_bit_slice_6541;
      p7_bit_slice_6542 <= p7_data_enable ? p6_bit_slice_6542 : p7_bit_slice_6542;
      p7_bit_slice_6543 <= p7_data_enable ? p6_bit_slice_6543 : p7_bit_slice_6543;
      p7_bit_slice_6544 <= p7_data_enable ? p6_bit_slice_6544 : p7_bit_slice_6544;
      p7_bit_slice_6545 <= p7_data_enable ? p6_bit_slice_6545 : p7_bit_slice_6545;
      p7_bit_slice_6546 <= p7_data_enable ? p6_bit_slice_6546 : p7_bit_slice_6546;
      p7_bit_slice_6547 <= p7_data_enable ? p6_bit_slice_6547 : p7_bit_slice_6547;
      p7_bit_slice_6548 <= p7_data_enable ? p6_bit_slice_6548 : p7_bit_slice_6548;
      p7_bit_slice_6549 <= p7_data_enable ? p6_bit_slice_6549 : p7_bit_slice_6549;
      p7_bit_slice_6550 <= p7_data_enable ? p6_bit_slice_6550 : p7_bit_slice_6550;
      p7_bit_slice_6551 <= p7_data_enable ? p6_bit_slice_6551 : p7_bit_slice_6551;
      p7_bit_slice_6552 <= p7_data_enable ? p6_bit_slice_6552 : p7_bit_slice_6552;
      p7_bit_slice_6553 <= p7_data_enable ? p6_bit_slice_6553 : p7_bit_slice_6553;
      p7_bit_slice_6554 <= p7_data_enable ? p6_bit_slice_6554 : p7_bit_slice_6554;
      p7_bit_slice_6555 <= p7_data_enable ? p6_bit_slice_6555 : p7_bit_slice_6555;
      p7_negated <= p7_data_enable ? p6_negated : p7_negated;
      p8_b <= p8_data_enable ? p7_b : p8_b;
      p8_uge_6629 <= p8_data_enable ? p7_uge_6629 : p8_uge_6629;
      p8_bivisor__1 <= p8_data_enable ? p7_bivisor__1 : p8_bivisor__1;
      p8_uge_6637 <= p8_data_enable ? p7_uge_6637 : p8_uge_6637;
      p8_uge_6719 <= p8_data_enable ? p7_uge_6719 : p8_uge_6719;
      p8_uge_6801 <= p8_data_enable ? p7_uge_6801 : p8_uge_6801;
      p8_uge_6881 <= p8_data_enable ? p7_uge_6881 : p8_uge_6881;
      p8_uge_6963 <= p8_data_enable ? p7_uge_6963 : p8_uge_6963;
      p8_uge_6969 <= p8_data_enable ? p7_uge_6969 : p8_uge_6969;
      p8_uge_7049 <= p8_data_enable ? p7_uge_7049 : p8_uge_7049;
      p8_uge_7131 <= p8_data_enable ? p7_uge_7131 : p8_uge_7131;
      p8_uge_7211 <= p8_data_enable ? uge_7211 : p8_uge_7211;
      p8_r__74 <= p8_data_enable ? r__74 : p8_r__74;
      p8_bit_slice_6534 <= p8_data_enable ? p7_bit_slice_6534 : p8_bit_slice_6534;
      p8_bit_slice_7214 <= p8_data_enable ? bit_slice_7214 : p8_bit_slice_7214;
      p8_bit_slice_6535 <= p8_data_enable ? p7_bit_slice_6535 : p8_bit_slice_6535;
      p8_bit_slice_6536 <= p8_data_enable ? p7_bit_slice_6536 : p8_bit_slice_6536;
      p8_bit_slice_6537 <= p8_data_enable ? p7_bit_slice_6537 : p8_bit_slice_6537;
      p8_bit_slice_6538 <= p8_data_enable ? p7_bit_slice_6538 : p8_bit_slice_6538;
      p8_bit_slice_6539 <= p8_data_enable ? p7_bit_slice_6539 : p8_bit_slice_6539;
      p8_bit_slice_6540 <= p8_data_enable ? p7_bit_slice_6540 : p8_bit_slice_6540;
      p8_bit_slice_6541 <= p8_data_enable ? p7_bit_slice_6541 : p8_bit_slice_6541;
      p8_bit_slice_6542 <= p8_data_enable ? p7_bit_slice_6542 : p8_bit_slice_6542;
      p8_bit_slice_6543 <= p8_data_enable ? p7_bit_slice_6543 : p8_bit_slice_6543;
      p8_bit_slice_6544 <= p8_data_enable ? p7_bit_slice_6544 : p8_bit_slice_6544;
      p8_bit_slice_6545 <= p8_data_enable ? p7_bit_slice_6545 : p8_bit_slice_6545;
      p8_bit_slice_6546 <= p8_data_enable ? p7_bit_slice_6546 : p8_bit_slice_6546;
      p8_bit_slice_6547 <= p8_data_enable ? p7_bit_slice_6547 : p8_bit_slice_6547;
      p8_bit_slice_6548 <= p8_data_enable ? p7_bit_slice_6548 : p8_bit_slice_6548;
      p8_bit_slice_6549 <= p8_data_enable ? p7_bit_slice_6549 : p8_bit_slice_6549;
      p8_bit_slice_6550 <= p8_data_enable ? p7_bit_slice_6550 : p8_bit_slice_6550;
      p8_bit_slice_6551 <= p8_data_enable ? p7_bit_slice_6551 : p8_bit_slice_6551;
      p8_bit_slice_6552 <= p8_data_enable ? p7_bit_slice_6552 : p8_bit_slice_6552;
      p8_bit_slice_6553 <= p8_data_enable ? p7_bit_slice_6553 : p8_bit_slice_6553;
      p8_bit_slice_6554 <= p8_data_enable ? p7_bit_slice_6554 : p8_bit_slice_6554;
      p8_bit_slice_6555 <= p8_data_enable ? p7_bit_slice_6555 : p8_bit_slice_6555;
      p8_negated <= p8_data_enable ? p7_negated : p8_negated;
      p9_b <= p9_data_enable ? p8_b : p9_b;
      p9_uge_6629 <= p9_data_enable ? p8_uge_6629 : p9_uge_6629;
      p9_bivisor__1 <= p9_data_enable ? p8_bivisor__1 : p9_bivisor__1;
      p9_uge_6637 <= p9_data_enable ? p8_uge_6637 : p9_uge_6637;
      p9_uge_6719 <= p9_data_enable ? p8_uge_6719 : p9_uge_6719;
      p9_uge_6801 <= p9_data_enable ? p8_uge_6801 : p9_uge_6801;
      p9_uge_6881 <= p9_data_enable ? p8_uge_6881 : p9_uge_6881;
      p9_uge_6963 <= p9_data_enable ? p8_uge_6963 : p9_uge_6963;
      p9_uge_6969 <= p9_data_enable ? p8_uge_6969 : p9_uge_6969;
      p9_uge_7049 <= p9_data_enable ? p8_uge_7049 : p9_uge_7049;
      p9_uge_7131 <= p9_data_enable ? p8_uge_7131 : p9_uge_7131;
      p9_uge_7211 <= p9_data_enable ? p8_uge_7211 : p9_uge_7211;
      p9_uge_7293 <= p9_data_enable ? uge_7293 : p9_uge_7293;
      p9_concat_7298 <= p9_data_enable ? concat_7298 : p9_concat_7298;
      p9_uge_7299 <= p9_data_enable ? uge_7299 : p9_uge_7299;
      p9_bit_slice_6536 <= p9_data_enable ? p8_bit_slice_6536 : p9_bit_slice_6536;
      p9_bit_slice_6537 <= p9_data_enable ? p8_bit_slice_6537 : p9_bit_slice_6537;
      p9_bit_slice_6538 <= p9_data_enable ? p8_bit_slice_6538 : p9_bit_slice_6538;
      p9_bit_slice_6539 <= p9_data_enable ? p8_bit_slice_6539 : p9_bit_slice_6539;
      p9_bit_slice_6540 <= p9_data_enable ? p8_bit_slice_6540 : p9_bit_slice_6540;
      p9_bit_slice_6541 <= p9_data_enable ? p8_bit_slice_6541 : p9_bit_slice_6541;
      p9_bit_slice_6542 <= p9_data_enable ? p8_bit_slice_6542 : p9_bit_slice_6542;
      p9_bit_slice_6543 <= p9_data_enable ? p8_bit_slice_6543 : p9_bit_slice_6543;
      p9_bit_slice_6544 <= p9_data_enable ? p8_bit_slice_6544 : p9_bit_slice_6544;
      p9_bit_slice_6545 <= p9_data_enable ? p8_bit_slice_6545 : p9_bit_slice_6545;
      p9_bit_slice_6546 <= p9_data_enable ? p8_bit_slice_6546 : p9_bit_slice_6546;
      p9_bit_slice_6547 <= p9_data_enable ? p8_bit_slice_6547 : p9_bit_slice_6547;
      p9_bit_slice_6548 <= p9_data_enable ? p8_bit_slice_6548 : p9_bit_slice_6548;
      p9_bit_slice_6549 <= p9_data_enable ? p8_bit_slice_6549 : p9_bit_slice_6549;
      p9_bit_slice_6550 <= p9_data_enable ? p8_bit_slice_6550 : p9_bit_slice_6550;
      p9_bit_slice_6551 <= p9_data_enable ? p8_bit_slice_6551 : p9_bit_slice_6551;
      p9_bit_slice_6552 <= p9_data_enable ? p8_bit_slice_6552 : p9_bit_slice_6552;
      p9_bit_slice_6553 <= p9_data_enable ? p8_bit_slice_6553 : p9_bit_slice_6553;
      p9_bit_slice_6554 <= p9_data_enable ? p8_bit_slice_6554 : p9_bit_slice_6554;
      p9_bit_slice_6555 <= p9_data_enable ? p8_bit_slice_6555 : p9_bit_slice_6555;
      p9_negated <= p9_data_enable ? p8_negated : p9_negated;
      p10_b <= p10_data_enable ? p9_b : p10_b;
      p10_uge_6629 <= p10_data_enable ? p9_uge_6629 : p10_uge_6629;
      p10_bivisor__1 <= p10_data_enable ? p9_bivisor__1 : p10_bivisor__1;
      p10_uge_6637 <= p10_data_enable ? p9_uge_6637 : p10_uge_6637;
      p10_uge_6719 <= p10_data_enable ? p9_uge_6719 : p10_uge_6719;
      p10_uge_6801 <= p10_data_enable ? p9_uge_6801 : p10_uge_6801;
      p10_uge_6881 <= p10_data_enable ? p9_uge_6881 : p10_uge_6881;
      p10_uge_6963 <= p10_data_enable ? p9_uge_6963 : p10_uge_6963;
      p10_uge_6969 <= p10_data_enable ? p9_uge_6969 : p10_uge_6969;
      p10_uge_7049 <= p10_data_enable ? p9_uge_7049 : p10_uge_7049;
      p10_uge_7131 <= p10_data_enable ? p9_uge_7131 : p10_uge_7131;
      p10_uge_7211 <= p10_data_enable ? p9_uge_7211 : p10_uge_7211;
      p10_uge_7293 <= p10_data_enable ? p9_uge_7293 : p10_uge_7293;
      p10_uge_7299 <= p10_data_enable ? p9_uge_7299 : p10_uge_7299;
      p10_concat_7378 <= p10_data_enable ? concat_7378 : p10_concat_7378;
      p10_uge_7379 <= p10_data_enable ? uge_7379 : p10_uge_7379;
      p10_sub_7380 <= p10_data_enable ? sub_7380 : p10_sub_7380;
      p10_bit_slice_6537 <= p10_data_enable ? p9_bit_slice_6537 : p10_bit_slice_6537;
      p10_bit_slice_6538 <= p10_data_enable ? p9_bit_slice_6538 : p10_bit_slice_6538;
      p10_bit_slice_6539 <= p10_data_enable ? p9_bit_slice_6539 : p10_bit_slice_6539;
      p10_bit_slice_6540 <= p10_data_enable ? p9_bit_slice_6540 : p10_bit_slice_6540;
      p10_bit_slice_6541 <= p10_data_enable ? p9_bit_slice_6541 : p10_bit_slice_6541;
      p10_bit_slice_6542 <= p10_data_enable ? p9_bit_slice_6542 : p10_bit_slice_6542;
      p10_bit_slice_6543 <= p10_data_enable ? p9_bit_slice_6543 : p10_bit_slice_6543;
      p10_bit_slice_6544 <= p10_data_enable ? p9_bit_slice_6544 : p10_bit_slice_6544;
      p10_bit_slice_6545 <= p10_data_enable ? p9_bit_slice_6545 : p10_bit_slice_6545;
      p10_bit_slice_6546 <= p10_data_enable ? p9_bit_slice_6546 : p10_bit_slice_6546;
      p10_bit_slice_6547 <= p10_data_enable ? p9_bit_slice_6547 : p10_bit_slice_6547;
      p10_bit_slice_6548 <= p10_data_enable ? p9_bit_slice_6548 : p10_bit_slice_6548;
      p10_bit_slice_6549 <= p10_data_enable ? p9_bit_slice_6549 : p10_bit_slice_6549;
      p10_bit_slice_6550 <= p10_data_enable ? p9_bit_slice_6550 : p10_bit_slice_6550;
      p10_bit_slice_6551 <= p10_data_enable ? p9_bit_slice_6551 : p10_bit_slice_6551;
      p10_bit_slice_6552 <= p10_data_enable ? p9_bit_slice_6552 : p10_bit_slice_6552;
      p10_bit_slice_6553 <= p10_data_enable ? p9_bit_slice_6553 : p10_bit_slice_6553;
      p10_bit_slice_6554 <= p10_data_enable ? p9_bit_slice_6554 : p10_bit_slice_6554;
      p10_bit_slice_6555 <= p10_data_enable ? p9_bit_slice_6555 : p10_bit_slice_6555;
      p10_negated <= p10_data_enable ? p9_negated : p10_negated;
      p11_b <= p11_data_enable ? p10_b : p11_b;
      p11_uge_6629 <= p11_data_enable ? p10_uge_6629 : p11_uge_6629;
      p11_bivisor__1 <= p11_data_enable ? p10_bivisor__1 : p11_bivisor__1;
      p11_uge_6637 <= p11_data_enable ? p10_uge_6637 : p11_uge_6637;
      p11_uge_6719 <= p11_data_enable ? p10_uge_6719 : p11_uge_6719;
      p11_uge_6801 <= p11_data_enable ? p10_uge_6801 : p11_uge_6801;
      p11_uge_6881 <= p11_data_enable ? p10_uge_6881 : p11_uge_6881;
      p11_uge_6963 <= p11_data_enable ? p10_uge_6963 : p11_uge_6963;
      p11_uge_6969 <= p11_data_enable ? p10_uge_6969 : p11_uge_6969;
      p11_uge_7049 <= p11_data_enable ? p10_uge_7049 : p11_uge_7049;
      p11_uge_7131 <= p11_data_enable ? p10_uge_7131 : p11_uge_7131;
      p11_uge_7211 <= p11_data_enable ? p10_uge_7211 : p11_uge_7211;
      p11_uge_7293 <= p11_data_enable ? p10_uge_7293 : p11_uge_7293;
      p11_uge_7299 <= p11_data_enable ? p10_uge_7299 : p11_uge_7299;
      p11_uge_7379 <= p11_data_enable ? p10_uge_7379 : p11_uge_7379;
      p11_uge_7461 <= p11_data_enable ? uge_7461 : p11_uge_7461;
      p11_r__78 <= p11_data_enable ? r__78 : p11_r__78;
      p11_bit_slice_6538 <= p11_data_enable ? p10_bit_slice_6538 : p11_bit_slice_6538;
      p11_bit_slice_6539 <= p11_data_enable ? p10_bit_slice_6539 : p11_bit_slice_6539;
      p11_bit_slice_6540 <= p11_data_enable ? p10_bit_slice_6540 : p11_bit_slice_6540;
      p11_bit_slice_6541 <= p11_data_enable ? p10_bit_slice_6541 : p11_bit_slice_6541;
      p11_bit_slice_6542 <= p11_data_enable ? p10_bit_slice_6542 : p11_bit_slice_6542;
      p11_bit_slice_6543 <= p11_data_enable ? p10_bit_slice_6543 : p11_bit_slice_6543;
      p11_bit_slice_6544 <= p11_data_enable ? p10_bit_slice_6544 : p11_bit_slice_6544;
      p11_bit_slice_6545 <= p11_data_enable ? p10_bit_slice_6545 : p11_bit_slice_6545;
      p11_bit_slice_6546 <= p11_data_enable ? p10_bit_slice_6546 : p11_bit_slice_6546;
      p11_bit_slice_6547 <= p11_data_enable ? p10_bit_slice_6547 : p11_bit_slice_6547;
      p11_bit_slice_6548 <= p11_data_enable ? p10_bit_slice_6548 : p11_bit_slice_6548;
      p11_bit_slice_6549 <= p11_data_enable ? p10_bit_slice_6549 : p11_bit_slice_6549;
      p11_bit_slice_6550 <= p11_data_enable ? p10_bit_slice_6550 : p11_bit_slice_6550;
      p11_bit_slice_6551 <= p11_data_enable ? p10_bit_slice_6551 : p11_bit_slice_6551;
      p11_bit_slice_6552 <= p11_data_enable ? p10_bit_slice_6552 : p11_bit_slice_6552;
      p11_bit_slice_6553 <= p11_data_enable ? p10_bit_slice_6553 : p11_bit_slice_6553;
      p11_bit_slice_6554 <= p11_data_enable ? p10_bit_slice_6554 : p11_bit_slice_6554;
      p11_bit_slice_6555 <= p11_data_enable ? p10_bit_slice_6555 : p11_bit_slice_6555;
      p11_negated <= p11_data_enable ? p10_negated : p11_negated;
      p12_b <= p12_data_enable ? p11_b : p12_b;
      p12_uge_6629 <= p12_data_enable ? p11_uge_6629 : p12_uge_6629;
      p12_bivisor__1 <= p12_data_enable ? p11_bivisor__1 : p12_bivisor__1;
      p12_uge_6637 <= p12_data_enable ? p11_uge_6637 : p12_uge_6637;
      p12_uge_6719 <= p12_data_enable ? p11_uge_6719 : p12_uge_6719;
      p12_uge_6801 <= p12_data_enable ? p11_uge_6801 : p12_uge_6801;
      p12_uge_6881 <= p12_data_enable ? p11_uge_6881 : p12_uge_6881;
      p12_uge_6963 <= p12_data_enable ? p11_uge_6963 : p12_uge_6963;
      p12_uge_6969 <= p12_data_enable ? p11_uge_6969 : p12_uge_6969;
      p12_uge_7049 <= p12_data_enable ? p11_uge_7049 : p12_uge_7049;
      p12_uge_7131 <= p12_data_enable ? p11_uge_7131 : p12_uge_7131;
      p12_uge_7211 <= p12_data_enable ? p11_uge_7211 : p12_uge_7211;
      p12_uge_7293 <= p12_data_enable ? p11_uge_7293 : p12_uge_7293;
      p12_uge_7299 <= p12_data_enable ? p11_uge_7299 : p12_uge_7299;
      p12_uge_7379 <= p12_data_enable ? p11_uge_7379 : p12_uge_7379;
      p12_uge_7461 <= p12_data_enable ? p11_uge_7461 : p12_uge_7461;
      p12_uge_7541 <= p12_data_enable ? uge_7541 : p12_uge_7541;
      p12_r__79 <= p12_data_enable ? r__79 : p12_r__79;
      p12_bit_slice_6539 <= p12_data_enable ? p11_bit_slice_6539 : p12_bit_slice_6539;
      p12_bit_slice_7544 <= p12_data_enable ? bit_slice_7544 : p12_bit_slice_7544;
      p12_bit_slice_6540 <= p12_data_enable ? p11_bit_slice_6540 : p12_bit_slice_6540;
      p12_bit_slice_6541 <= p12_data_enable ? p11_bit_slice_6541 : p12_bit_slice_6541;
      p12_bit_slice_6542 <= p12_data_enable ? p11_bit_slice_6542 : p12_bit_slice_6542;
      p12_bit_slice_6543 <= p12_data_enable ? p11_bit_slice_6543 : p12_bit_slice_6543;
      p12_bit_slice_6544 <= p12_data_enable ? p11_bit_slice_6544 : p12_bit_slice_6544;
      p12_bit_slice_6545 <= p12_data_enable ? p11_bit_slice_6545 : p12_bit_slice_6545;
      p12_bit_slice_6546 <= p12_data_enable ? p11_bit_slice_6546 : p12_bit_slice_6546;
      p12_bit_slice_6547 <= p12_data_enable ? p11_bit_slice_6547 : p12_bit_slice_6547;
      p12_bit_slice_6548 <= p12_data_enable ? p11_bit_slice_6548 : p12_bit_slice_6548;
      p12_bit_slice_6549 <= p12_data_enable ? p11_bit_slice_6549 : p12_bit_slice_6549;
      p12_bit_slice_6550 <= p12_data_enable ? p11_bit_slice_6550 : p12_bit_slice_6550;
      p12_bit_slice_6551 <= p12_data_enable ? p11_bit_slice_6551 : p12_bit_slice_6551;
      p12_bit_slice_6552 <= p12_data_enable ? p11_bit_slice_6552 : p12_bit_slice_6552;
      p12_bit_slice_6553 <= p12_data_enable ? p11_bit_slice_6553 : p12_bit_slice_6553;
      p12_bit_slice_6554 <= p12_data_enable ? p11_bit_slice_6554 : p12_bit_slice_6554;
      p12_bit_slice_6555 <= p12_data_enable ? p11_bit_slice_6555 : p12_bit_slice_6555;
      p12_negated <= p12_data_enable ? p11_negated : p12_negated;
      p13_b <= p13_data_enable ? p12_b : p13_b;
      p13_uge_6629 <= p13_data_enable ? p12_uge_6629 : p13_uge_6629;
      p13_bivisor__1 <= p13_data_enable ? p12_bivisor__1 : p13_bivisor__1;
      p13_uge_6637 <= p13_data_enable ? p12_uge_6637 : p13_uge_6637;
      p13_uge_6719 <= p13_data_enable ? p12_uge_6719 : p13_uge_6719;
      p13_uge_6801 <= p13_data_enable ? p12_uge_6801 : p13_uge_6801;
      p13_uge_6881 <= p13_data_enable ? p12_uge_6881 : p13_uge_6881;
      p13_uge_6963 <= p13_data_enable ? p12_uge_6963 : p13_uge_6963;
      p13_uge_6969 <= p13_data_enable ? p12_uge_6969 : p13_uge_6969;
      p13_uge_7049 <= p13_data_enable ? p12_uge_7049 : p13_uge_7049;
      p13_uge_7131 <= p13_data_enable ? p12_uge_7131 : p13_uge_7131;
      p13_uge_7211 <= p13_data_enable ? p12_uge_7211 : p13_uge_7211;
      p13_uge_7293 <= p13_data_enable ? p12_uge_7293 : p13_uge_7293;
      p13_uge_7299 <= p13_data_enable ? p12_uge_7299 : p13_uge_7299;
      p13_uge_7379 <= p13_data_enable ? p12_uge_7379 : p13_uge_7379;
      p13_uge_7461 <= p13_data_enable ? p12_uge_7461 : p13_uge_7461;
      p13_uge_7541 <= p13_data_enable ? p12_uge_7541 : p13_uge_7541;
      p13_uge_7623 <= p13_data_enable ? uge_7623 : p13_uge_7623;
      p13_concat_7628 <= p13_data_enable ? concat_7628 : p13_concat_7628;
      p13_uge_7629 <= p13_data_enable ? uge_7629 : p13_uge_7629;
      p13_bit_slice_6541 <= p13_data_enable ? p12_bit_slice_6541 : p13_bit_slice_6541;
      p13_bit_slice_6542 <= p13_data_enable ? p12_bit_slice_6542 : p13_bit_slice_6542;
      p13_bit_slice_6543 <= p13_data_enable ? p12_bit_slice_6543 : p13_bit_slice_6543;
      p13_bit_slice_6544 <= p13_data_enable ? p12_bit_slice_6544 : p13_bit_slice_6544;
      p13_bit_slice_6545 <= p13_data_enable ? p12_bit_slice_6545 : p13_bit_slice_6545;
      p13_bit_slice_6546 <= p13_data_enable ? p12_bit_slice_6546 : p13_bit_slice_6546;
      p13_bit_slice_6547 <= p13_data_enable ? p12_bit_slice_6547 : p13_bit_slice_6547;
      p13_bit_slice_6548 <= p13_data_enable ? p12_bit_slice_6548 : p13_bit_slice_6548;
      p13_bit_slice_6549 <= p13_data_enable ? p12_bit_slice_6549 : p13_bit_slice_6549;
      p13_bit_slice_6550 <= p13_data_enable ? p12_bit_slice_6550 : p13_bit_slice_6550;
      p13_bit_slice_6551 <= p13_data_enable ? p12_bit_slice_6551 : p13_bit_slice_6551;
      p13_bit_slice_6552 <= p13_data_enable ? p12_bit_slice_6552 : p13_bit_slice_6552;
      p13_bit_slice_6553 <= p13_data_enable ? p12_bit_slice_6553 : p13_bit_slice_6553;
      p13_bit_slice_6554 <= p13_data_enable ? p12_bit_slice_6554 : p13_bit_slice_6554;
      p13_bit_slice_6555 <= p13_data_enable ? p12_bit_slice_6555 : p13_bit_slice_6555;
      p13_negated <= p13_data_enable ? p12_negated : p13_negated;
      p14_b <= p14_data_enable ? p13_b : p14_b;
      p14_uge_6629 <= p14_data_enable ? p13_uge_6629 : p14_uge_6629;
      p14_bivisor__1 <= p14_data_enable ? p13_bivisor__1 : p14_bivisor__1;
      p14_uge_6637 <= p14_data_enable ? p13_uge_6637 : p14_uge_6637;
      p14_uge_6719 <= p14_data_enable ? p13_uge_6719 : p14_uge_6719;
      p14_uge_6801 <= p14_data_enable ? p13_uge_6801 : p14_uge_6801;
      p14_uge_6881 <= p14_data_enable ? p13_uge_6881 : p14_uge_6881;
      p14_uge_6963 <= p14_data_enable ? p13_uge_6963 : p14_uge_6963;
      p14_uge_6969 <= p14_data_enable ? p13_uge_6969 : p14_uge_6969;
      p14_uge_7049 <= p14_data_enable ? p13_uge_7049 : p14_uge_7049;
      p14_uge_7131 <= p14_data_enable ? p13_uge_7131 : p14_uge_7131;
      p14_uge_7211 <= p14_data_enable ? p13_uge_7211 : p14_uge_7211;
      p14_uge_7293 <= p14_data_enable ? p13_uge_7293 : p14_uge_7293;
      p14_uge_7299 <= p14_data_enable ? p13_uge_7299 : p14_uge_7299;
      p14_uge_7379 <= p14_data_enable ? p13_uge_7379 : p14_uge_7379;
      p14_uge_7461 <= p14_data_enable ? p13_uge_7461 : p14_uge_7461;
      p14_uge_7541 <= p14_data_enable ? p13_uge_7541 : p14_uge_7541;
      p14_uge_7623 <= p14_data_enable ? p13_uge_7623 : p14_uge_7623;
      p14_uge_7629 <= p14_data_enable ? p13_uge_7629 : p14_uge_7629;
      p14_concat_7708 <= p14_data_enable ? concat_7708 : p14_concat_7708;
      p14_uge_7709 <= p14_data_enable ? uge_7709 : p14_uge_7709;
      p14_sub_7710 <= p14_data_enable ? sub_7710 : p14_sub_7710;
      p14_bit_slice_6542 <= p14_data_enable ? p13_bit_slice_6542 : p14_bit_slice_6542;
      p14_bit_slice_6543 <= p14_data_enable ? p13_bit_slice_6543 : p14_bit_slice_6543;
      p14_bit_slice_6544 <= p14_data_enable ? p13_bit_slice_6544 : p14_bit_slice_6544;
      p14_bit_slice_6545 <= p14_data_enable ? p13_bit_slice_6545 : p14_bit_slice_6545;
      p14_bit_slice_6546 <= p14_data_enable ? p13_bit_slice_6546 : p14_bit_slice_6546;
      p14_bit_slice_6547 <= p14_data_enable ? p13_bit_slice_6547 : p14_bit_slice_6547;
      p14_bit_slice_6548 <= p14_data_enable ? p13_bit_slice_6548 : p14_bit_slice_6548;
      p14_bit_slice_6549 <= p14_data_enable ? p13_bit_slice_6549 : p14_bit_slice_6549;
      p14_bit_slice_6550 <= p14_data_enable ? p13_bit_slice_6550 : p14_bit_slice_6550;
      p14_bit_slice_6551 <= p14_data_enable ? p13_bit_slice_6551 : p14_bit_slice_6551;
      p14_bit_slice_6552 <= p14_data_enable ? p13_bit_slice_6552 : p14_bit_slice_6552;
      p14_bit_slice_6553 <= p14_data_enable ? p13_bit_slice_6553 : p14_bit_slice_6553;
      p14_bit_slice_6554 <= p14_data_enable ? p13_bit_slice_6554 : p14_bit_slice_6554;
      p14_bit_slice_6555 <= p14_data_enable ? p13_bit_slice_6555 : p14_bit_slice_6555;
      p14_negated <= p14_data_enable ? p13_negated : p14_negated;
      p15_b <= p15_data_enable ? p14_b : p15_b;
      p15_uge_6629 <= p15_data_enable ? p14_uge_6629 : p15_uge_6629;
      p15_bivisor__1 <= p15_data_enable ? p14_bivisor__1 : p15_bivisor__1;
      p15_uge_6637 <= p15_data_enable ? p14_uge_6637 : p15_uge_6637;
      p15_uge_6719 <= p15_data_enable ? p14_uge_6719 : p15_uge_6719;
      p15_uge_6801 <= p15_data_enable ? p14_uge_6801 : p15_uge_6801;
      p15_uge_6881 <= p15_data_enable ? p14_uge_6881 : p15_uge_6881;
      p15_uge_6963 <= p15_data_enable ? p14_uge_6963 : p15_uge_6963;
      p15_uge_6969 <= p15_data_enable ? p14_uge_6969 : p15_uge_6969;
      p15_uge_7049 <= p15_data_enable ? p14_uge_7049 : p15_uge_7049;
      p15_uge_7131 <= p15_data_enable ? p14_uge_7131 : p15_uge_7131;
      p15_uge_7211 <= p15_data_enable ? p14_uge_7211 : p15_uge_7211;
      p15_uge_7293 <= p15_data_enable ? p14_uge_7293 : p15_uge_7293;
      p15_uge_7299 <= p15_data_enable ? p14_uge_7299 : p15_uge_7299;
      p15_uge_7379 <= p15_data_enable ? p14_uge_7379 : p15_uge_7379;
      p15_uge_7461 <= p15_data_enable ? p14_uge_7461 : p15_uge_7461;
      p15_uge_7541 <= p15_data_enable ? p14_uge_7541 : p15_uge_7541;
      p15_uge_7623 <= p15_data_enable ? p14_uge_7623 : p15_uge_7623;
      p15_uge_7629 <= p15_data_enable ? p14_uge_7629 : p15_uge_7629;
      p15_uge_7709 <= p15_data_enable ? p14_uge_7709 : p15_uge_7709;
      p15_uge_7791 <= p15_data_enable ? uge_7791 : p15_uge_7791;
      p15_r__83 <= p15_data_enable ? r__83 : p15_r__83;
      p15_bit_slice_6543 <= p15_data_enable ? p14_bit_slice_6543 : p15_bit_slice_6543;
      p15_bit_slice_6544 <= p15_data_enable ? p14_bit_slice_6544 : p15_bit_slice_6544;
      p15_bit_slice_6545 <= p15_data_enable ? p14_bit_slice_6545 : p15_bit_slice_6545;
      p15_bit_slice_6546 <= p15_data_enable ? p14_bit_slice_6546 : p15_bit_slice_6546;
      p15_bit_slice_6547 <= p15_data_enable ? p14_bit_slice_6547 : p15_bit_slice_6547;
      p15_bit_slice_6548 <= p15_data_enable ? p14_bit_slice_6548 : p15_bit_slice_6548;
      p15_bit_slice_6549 <= p15_data_enable ? p14_bit_slice_6549 : p15_bit_slice_6549;
      p15_bit_slice_6550 <= p15_data_enable ? p14_bit_slice_6550 : p15_bit_slice_6550;
      p15_bit_slice_6551 <= p15_data_enable ? p14_bit_slice_6551 : p15_bit_slice_6551;
      p15_bit_slice_6552 <= p15_data_enable ? p14_bit_slice_6552 : p15_bit_slice_6552;
      p15_bit_slice_6553 <= p15_data_enable ? p14_bit_slice_6553 : p15_bit_slice_6553;
      p15_bit_slice_6554 <= p15_data_enable ? p14_bit_slice_6554 : p15_bit_slice_6554;
      p15_bit_slice_6555 <= p15_data_enable ? p14_bit_slice_6555 : p15_bit_slice_6555;
      p15_negated <= p15_data_enable ? p14_negated : p15_negated;
      p16_b <= p16_data_enable ? p15_b : p16_b;
      p16_uge_6629 <= p16_data_enable ? p15_uge_6629 : p16_uge_6629;
      p16_bivisor__1 <= p16_data_enable ? p15_bivisor__1 : p16_bivisor__1;
      p16_uge_6637 <= p16_data_enable ? p15_uge_6637 : p16_uge_6637;
      p16_uge_6719 <= p16_data_enable ? p15_uge_6719 : p16_uge_6719;
      p16_uge_6801 <= p16_data_enable ? p15_uge_6801 : p16_uge_6801;
      p16_uge_6881 <= p16_data_enable ? p15_uge_6881 : p16_uge_6881;
      p16_uge_6963 <= p16_data_enable ? p15_uge_6963 : p16_uge_6963;
      p16_uge_6969 <= p16_data_enable ? p15_uge_6969 : p16_uge_6969;
      p16_uge_7049 <= p16_data_enable ? p15_uge_7049 : p16_uge_7049;
      p16_uge_7131 <= p16_data_enable ? p15_uge_7131 : p16_uge_7131;
      p16_uge_7211 <= p16_data_enable ? p15_uge_7211 : p16_uge_7211;
      p16_uge_7293 <= p16_data_enable ? p15_uge_7293 : p16_uge_7293;
      p16_uge_7299 <= p16_data_enable ? p15_uge_7299 : p16_uge_7299;
      p16_uge_7379 <= p16_data_enable ? p15_uge_7379 : p16_uge_7379;
      p16_uge_7461 <= p16_data_enable ? p15_uge_7461 : p16_uge_7461;
      p16_uge_7541 <= p16_data_enable ? p15_uge_7541 : p16_uge_7541;
      p16_uge_7623 <= p16_data_enable ? p15_uge_7623 : p16_uge_7623;
      p16_uge_7629 <= p16_data_enable ? p15_uge_7629 : p16_uge_7629;
      p16_uge_7709 <= p16_data_enable ? p15_uge_7709 : p16_uge_7709;
      p16_uge_7791 <= p16_data_enable ? p15_uge_7791 : p16_uge_7791;
      p16_uge_7871 <= p16_data_enable ? uge_7871 : p16_uge_7871;
      p16_r__84 <= p16_data_enable ? r__84 : p16_r__84;
      p16_bit_slice_6544 <= p16_data_enable ? p15_bit_slice_6544 : p16_bit_slice_6544;
      p16_bit_slice_7874 <= p16_data_enable ? bit_slice_7874 : p16_bit_slice_7874;
      p16_bit_slice_6545 <= p16_data_enable ? p15_bit_slice_6545 : p16_bit_slice_6545;
      p16_bit_slice_6546 <= p16_data_enable ? p15_bit_slice_6546 : p16_bit_slice_6546;
      p16_bit_slice_6547 <= p16_data_enable ? p15_bit_slice_6547 : p16_bit_slice_6547;
      p16_bit_slice_6548 <= p16_data_enable ? p15_bit_slice_6548 : p16_bit_slice_6548;
      p16_bit_slice_6549 <= p16_data_enable ? p15_bit_slice_6549 : p16_bit_slice_6549;
      p16_bit_slice_6550 <= p16_data_enable ? p15_bit_slice_6550 : p16_bit_slice_6550;
      p16_bit_slice_6551 <= p16_data_enable ? p15_bit_slice_6551 : p16_bit_slice_6551;
      p16_bit_slice_6552 <= p16_data_enable ? p15_bit_slice_6552 : p16_bit_slice_6552;
      p16_bit_slice_6553 <= p16_data_enable ? p15_bit_slice_6553 : p16_bit_slice_6553;
      p16_bit_slice_6554 <= p16_data_enable ? p15_bit_slice_6554 : p16_bit_slice_6554;
      p16_bit_slice_6555 <= p16_data_enable ? p15_bit_slice_6555 : p16_bit_slice_6555;
      p16_negated <= p16_data_enable ? p15_negated : p16_negated;
      p17_b <= p17_data_enable ? p16_b : p17_b;
      p17_uge_6629 <= p17_data_enable ? p16_uge_6629 : p17_uge_6629;
      p17_bivisor__1 <= p17_data_enable ? p16_bivisor__1 : p17_bivisor__1;
      p17_uge_6637 <= p17_data_enable ? p16_uge_6637 : p17_uge_6637;
      p17_uge_6719 <= p17_data_enable ? p16_uge_6719 : p17_uge_6719;
      p17_uge_6801 <= p17_data_enable ? p16_uge_6801 : p17_uge_6801;
      p17_uge_6881 <= p17_data_enable ? p16_uge_6881 : p17_uge_6881;
      p17_uge_6963 <= p17_data_enable ? p16_uge_6963 : p17_uge_6963;
      p17_uge_6969 <= p17_data_enable ? p16_uge_6969 : p17_uge_6969;
      p17_uge_7049 <= p17_data_enable ? p16_uge_7049 : p17_uge_7049;
      p17_uge_7131 <= p17_data_enable ? p16_uge_7131 : p17_uge_7131;
      p17_uge_7211 <= p17_data_enable ? p16_uge_7211 : p17_uge_7211;
      p17_uge_7293 <= p17_data_enable ? p16_uge_7293 : p17_uge_7293;
      p17_uge_7299 <= p17_data_enable ? p16_uge_7299 : p17_uge_7299;
      p17_uge_7379 <= p17_data_enable ? p16_uge_7379 : p17_uge_7379;
      p17_uge_7461 <= p17_data_enable ? p16_uge_7461 : p17_uge_7461;
      p17_uge_7541 <= p17_data_enable ? p16_uge_7541 : p17_uge_7541;
      p17_uge_7623 <= p17_data_enable ? p16_uge_7623 : p17_uge_7623;
      p17_uge_7629 <= p17_data_enable ? p16_uge_7629 : p17_uge_7629;
      p17_uge_7709 <= p17_data_enable ? p16_uge_7709 : p17_uge_7709;
      p17_uge_7791 <= p17_data_enable ? p16_uge_7791 : p17_uge_7791;
      p17_uge_7871 <= p17_data_enable ? p16_uge_7871 : p17_uge_7871;
      p17_uge_7953 <= p17_data_enable ? uge_7953 : p17_uge_7953;
      p17_concat_7958 <= p17_data_enable ? concat_7958 : p17_concat_7958;
      p17_uge_7959 <= p17_data_enable ? uge_7959 : p17_uge_7959;
      p17_bit_slice_6546 <= p17_data_enable ? p16_bit_slice_6546 : p17_bit_slice_6546;
      p17_bit_slice_6547 <= p17_data_enable ? p16_bit_slice_6547 : p17_bit_slice_6547;
      p17_bit_slice_6548 <= p17_data_enable ? p16_bit_slice_6548 : p17_bit_slice_6548;
      p17_bit_slice_6549 <= p17_data_enable ? p16_bit_slice_6549 : p17_bit_slice_6549;
      p17_bit_slice_6550 <= p17_data_enable ? p16_bit_slice_6550 : p17_bit_slice_6550;
      p17_bit_slice_6551 <= p17_data_enable ? p16_bit_slice_6551 : p17_bit_slice_6551;
      p17_bit_slice_6552 <= p17_data_enable ? p16_bit_slice_6552 : p17_bit_slice_6552;
      p17_bit_slice_6553 <= p17_data_enable ? p16_bit_slice_6553 : p17_bit_slice_6553;
      p17_bit_slice_6554 <= p17_data_enable ? p16_bit_slice_6554 : p17_bit_slice_6554;
      p17_bit_slice_6555 <= p17_data_enable ? p16_bit_slice_6555 : p17_bit_slice_6555;
      p17_negated <= p17_data_enable ? p16_negated : p17_negated;
      p18_b <= p18_data_enable ? p17_b : p18_b;
      p18_uge_6629 <= p18_data_enable ? p17_uge_6629 : p18_uge_6629;
      p18_bivisor__1 <= p18_data_enable ? p17_bivisor__1 : p18_bivisor__1;
      p18_uge_6637 <= p18_data_enable ? p17_uge_6637 : p18_uge_6637;
      p18_uge_6719 <= p18_data_enable ? p17_uge_6719 : p18_uge_6719;
      p18_uge_6801 <= p18_data_enable ? p17_uge_6801 : p18_uge_6801;
      p18_uge_6881 <= p18_data_enable ? p17_uge_6881 : p18_uge_6881;
      p18_uge_6963 <= p18_data_enable ? p17_uge_6963 : p18_uge_6963;
      p18_uge_6969 <= p18_data_enable ? p17_uge_6969 : p18_uge_6969;
      p18_uge_7049 <= p18_data_enable ? p17_uge_7049 : p18_uge_7049;
      p18_uge_7131 <= p18_data_enable ? p17_uge_7131 : p18_uge_7131;
      p18_uge_7211 <= p18_data_enable ? p17_uge_7211 : p18_uge_7211;
      p18_uge_7293 <= p18_data_enable ? p17_uge_7293 : p18_uge_7293;
      p18_uge_7299 <= p18_data_enable ? p17_uge_7299 : p18_uge_7299;
      p18_uge_7379 <= p18_data_enable ? p17_uge_7379 : p18_uge_7379;
      p18_uge_7461 <= p18_data_enable ? p17_uge_7461 : p18_uge_7461;
      p18_uge_7541 <= p18_data_enable ? p17_uge_7541 : p18_uge_7541;
      p18_uge_7623 <= p18_data_enable ? p17_uge_7623 : p18_uge_7623;
      p18_uge_7629 <= p18_data_enable ? p17_uge_7629 : p18_uge_7629;
      p18_uge_7709 <= p18_data_enable ? p17_uge_7709 : p18_uge_7709;
      p18_uge_7791 <= p18_data_enable ? p17_uge_7791 : p18_uge_7791;
      p18_uge_7871 <= p18_data_enable ? p17_uge_7871 : p18_uge_7871;
      p18_uge_7953 <= p18_data_enable ? p17_uge_7953 : p18_uge_7953;
      p18_uge_7959 <= p18_data_enable ? p17_uge_7959 : p18_uge_7959;
      p18_concat_8038 <= p18_data_enable ? concat_8038 : p18_concat_8038;
      p18_uge_8039 <= p18_data_enable ? uge_8039 : p18_uge_8039;
      p18_sub_8040 <= p18_data_enable ? sub_8040 : p18_sub_8040;
      p18_bit_slice_6547 <= p18_data_enable ? p17_bit_slice_6547 : p18_bit_slice_6547;
      p18_bit_slice_6548 <= p18_data_enable ? p17_bit_slice_6548 : p18_bit_slice_6548;
      p18_bit_slice_6549 <= p18_data_enable ? p17_bit_slice_6549 : p18_bit_slice_6549;
      p18_bit_slice_6550 <= p18_data_enable ? p17_bit_slice_6550 : p18_bit_slice_6550;
      p18_bit_slice_6551 <= p18_data_enable ? p17_bit_slice_6551 : p18_bit_slice_6551;
      p18_bit_slice_6552 <= p18_data_enable ? p17_bit_slice_6552 : p18_bit_slice_6552;
      p18_bit_slice_6553 <= p18_data_enable ? p17_bit_slice_6553 : p18_bit_slice_6553;
      p18_bit_slice_6554 <= p18_data_enable ? p17_bit_slice_6554 : p18_bit_slice_6554;
      p18_bit_slice_6555 <= p18_data_enable ? p17_bit_slice_6555 : p18_bit_slice_6555;
      p18_negated <= p18_data_enable ? p17_negated : p18_negated;
      p19_b <= p19_data_enable ? p18_b : p19_b;
      p19_uge_6629 <= p19_data_enable ? p18_uge_6629 : p19_uge_6629;
      p19_bivisor__1 <= p19_data_enable ? p18_bivisor__1 : p19_bivisor__1;
      p19_uge_6637 <= p19_data_enable ? p18_uge_6637 : p19_uge_6637;
      p19_uge_6719 <= p19_data_enable ? p18_uge_6719 : p19_uge_6719;
      p19_uge_6801 <= p19_data_enable ? p18_uge_6801 : p19_uge_6801;
      p19_uge_6881 <= p19_data_enable ? p18_uge_6881 : p19_uge_6881;
      p19_uge_6963 <= p19_data_enable ? p18_uge_6963 : p19_uge_6963;
      p19_uge_6969 <= p19_data_enable ? p18_uge_6969 : p19_uge_6969;
      p19_uge_7049 <= p19_data_enable ? p18_uge_7049 : p19_uge_7049;
      p19_uge_7131 <= p19_data_enable ? p18_uge_7131 : p19_uge_7131;
      p19_uge_7211 <= p19_data_enable ? p18_uge_7211 : p19_uge_7211;
      p19_uge_7293 <= p19_data_enable ? p18_uge_7293 : p19_uge_7293;
      p19_uge_7299 <= p19_data_enable ? p18_uge_7299 : p19_uge_7299;
      p19_uge_7379 <= p19_data_enable ? p18_uge_7379 : p19_uge_7379;
      p19_uge_7461 <= p19_data_enable ? p18_uge_7461 : p19_uge_7461;
      p19_uge_7541 <= p19_data_enable ? p18_uge_7541 : p19_uge_7541;
      p19_uge_7623 <= p19_data_enable ? p18_uge_7623 : p19_uge_7623;
      p19_uge_7629 <= p19_data_enable ? p18_uge_7629 : p19_uge_7629;
      p19_uge_7709 <= p19_data_enable ? p18_uge_7709 : p19_uge_7709;
      p19_uge_7791 <= p19_data_enable ? p18_uge_7791 : p19_uge_7791;
      p19_uge_7871 <= p19_data_enable ? p18_uge_7871 : p19_uge_7871;
      p19_uge_7953 <= p19_data_enable ? p18_uge_7953 : p19_uge_7953;
      p19_uge_7959 <= p19_data_enable ? p18_uge_7959 : p19_uge_7959;
      p19_uge_8039 <= p19_data_enable ? p18_uge_8039 : p19_uge_8039;
      p19_uge_8121 <= p19_data_enable ? uge_8121 : p19_uge_8121;
      p19_r__88 <= p19_data_enable ? r__88 : p19_r__88;
      p19_bit_slice_6548 <= p19_data_enable ? p18_bit_slice_6548 : p19_bit_slice_6548;
      p19_bit_slice_6549 <= p19_data_enable ? p18_bit_slice_6549 : p19_bit_slice_6549;
      p19_bit_slice_6550 <= p19_data_enable ? p18_bit_slice_6550 : p19_bit_slice_6550;
      p19_bit_slice_6551 <= p19_data_enable ? p18_bit_slice_6551 : p19_bit_slice_6551;
      p19_bit_slice_6552 <= p19_data_enable ? p18_bit_slice_6552 : p19_bit_slice_6552;
      p19_bit_slice_6553 <= p19_data_enable ? p18_bit_slice_6553 : p19_bit_slice_6553;
      p19_bit_slice_6554 <= p19_data_enable ? p18_bit_slice_6554 : p19_bit_slice_6554;
      p19_bit_slice_6555 <= p19_data_enable ? p18_bit_slice_6555 : p19_bit_slice_6555;
      p19_negated <= p19_data_enable ? p18_negated : p19_negated;
      p20_b <= p20_data_enable ? p19_b : p20_b;
      p20_uge_6629 <= p20_data_enable ? p19_uge_6629 : p20_uge_6629;
      p20_bivisor__1 <= p20_data_enable ? p19_bivisor__1 : p20_bivisor__1;
      p20_uge_6637 <= p20_data_enable ? p19_uge_6637 : p20_uge_6637;
      p20_uge_6719 <= p20_data_enable ? p19_uge_6719 : p20_uge_6719;
      p20_uge_6801 <= p20_data_enable ? p19_uge_6801 : p20_uge_6801;
      p20_uge_6881 <= p20_data_enable ? p19_uge_6881 : p20_uge_6881;
      p20_uge_6963 <= p20_data_enable ? p19_uge_6963 : p20_uge_6963;
      p20_uge_6969 <= p20_data_enable ? p19_uge_6969 : p20_uge_6969;
      p20_uge_7049 <= p20_data_enable ? p19_uge_7049 : p20_uge_7049;
      p20_uge_7131 <= p20_data_enable ? p19_uge_7131 : p20_uge_7131;
      p20_uge_7211 <= p20_data_enable ? p19_uge_7211 : p20_uge_7211;
      p20_uge_7293 <= p20_data_enable ? p19_uge_7293 : p20_uge_7293;
      p20_uge_7299 <= p20_data_enable ? p19_uge_7299 : p20_uge_7299;
      p20_uge_7379 <= p20_data_enable ? p19_uge_7379 : p20_uge_7379;
      p20_uge_7461 <= p20_data_enable ? p19_uge_7461 : p20_uge_7461;
      p20_uge_7541 <= p20_data_enable ? p19_uge_7541 : p20_uge_7541;
      p20_uge_7623 <= p20_data_enable ? p19_uge_7623 : p20_uge_7623;
      p20_uge_7629 <= p20_data_enable ? p19_uge_7629 : p20_uge_7629;
      p20_uge_7709 <= p20_data_enable ? p19_uge_7709 : p20_uge_7709;
      p20_uge_7791 <= p20_data_enable ? p19_uge_7791 : p20_uge_7791;
      p20_uge_7871 <= p20_data_enable ? p19_uge_7871 : p20_uge_7871;
      p20_uge_7953 <= p20_data_enable ? p19_uge_7953 : p20_uge_7953;
      p20_uge_7959 <= p20_data_enable ? p19_uge_7959 : p20_uge_7959;
      p20_uge_8039 <= p20_data_enable ? p19_uge_8039 : p20_uge_8039;
      p20_uge_8121 <= p20_data_enable ? p19_uge_8121 : p20_uge_8121;
      p20_uge_8201 <= p20_data_enable ? uge_8201 : p20_uge_8201;
      p20_r__89 <= p20_data_enable ? r__89 : p20_r__89;
      p20_bit_slice_6549 <= p20_data_enable ? p19_bit_slice_6549 : p20_bit_slice_6549;
      p20_bit_slice_8204 <= p20_data_enable ? bit_slice_8204 : p20_bit_slice_8204;
      p20_bit_slice_6550 <= p20_data_enable ? p19_bit_slice_6550 : p20_bit_slice_6550;
      p20_bit_slice_6551 <= p20_data_enable ? p19_bit_slice_6551 : p20_bit_slice_6551;
      p20_bit_slice_6552 <= p20_data_enable ? p19_bit_slice_6552 : p20_bit_slice_6552;
      p20_bit_slice_6553 <= p20_data_enable ? p19_bit_slice_6553 : p20_bit_slice_6553;
      p20_bit_slice_6554 <= p20_data_enable ? p19_bit_slice_6554 : p20_bit_slice_6554;
      p20_bit_slice_6555 <= p20_data_enable ? p19_bit_slice_6555 : p20_bit_slice_6555;
      p20_negated <= p20_data_enable ? p19_negated : p20_negated;
      p21_b <= p21_data_enable ? p20_b : p21_b;
      p21_uge_6629 <= p21_data_enable ? p20_uge_6629 : p21_uge_6629;
      p21_bivisor__1 <= p21_data_enable ? p20_bivisor__1 : p21_bivisor__1;
      p21_uge_6637 <= p21_data_enable ? p20_uge_6637 : p21_uge_6637;
      p21_uge_6719 <= p21_data_enable ? p20_uge_6719 : p21_uge_6719;
      p21_uge_6801 <= p21_data_enable ? p20_uge_6801 : p21_uge_6801;
      p21_uge_6881 <= p21_data_enable ? p20_uge_6881 : p21_uge_6881;
      p21_uge_6963 <= p21_data_enable ? p20_uge_6963 : p21_uge_6963;
      p21_uge_6969 <= p21_data_enable ? p20_uge_6969 : p21_uge_6969;
      p21_uge_7049 <= p21_data_enable ? p20_uge_7049 : p21_uge_7049;
      p21_uge_7131 <= p21_data_enable ? p20_uge_7131 : p21_uge_7131;
      p21_uge_7211 <= p21_data_enable ? p20_uge_7211 : p21_uge_7211;
      p21_uge_7293 <= p21_data_enable ? p20_uge_7293 : p21_uge_7293;
      p21_uge_7299 <= p21_data_enable ? p20_uge_7299 : p21_uge_7299;
      p21_uge_7379 <= p21_data_enable ? p20_uge_7379 : p21_uge_7379;
      p21_uge_7461 <= p21_data_enable ? p20_uge_7461 : p21_uge_7461;
      p21_uge_7541 <= p21_data_enable ? p20_uge_7541 : p21_uge_7541;
      p21_uge_7623 <= p21_data_enable ? p20_uge_7623 : p21_uge_7623;
      p21_uge_7629 <= p21_data_enable ? p20_uge_7629 : p21_uge_7629;
      p21_uge_7709 <= p21_data_enable ? p20_uge_7709 : p21_uge_7709;
      p21_uge_7791 <= p21_data_enable ? p20_uge_7791 : p21_uge_7791;
      p21_uge_7871 <= p21_data_enable ? p20_uge_7871 : p21_uge_7871;
      p21_uge_7953 <= p21_data_enable ? p20_uge_7953 : p21_uge_7953;
      p21_uge_7959 <= p21_data_enable ? p20_uge_7959 : p21_uge_7959;
      p21_uge_8039 <= p21_data_enable ? p20_uge_8039 : p21_uge_8039;
      p21_uge_8121 <= p21_data_enable ? p20_uge_8121 : p21_uge_8121;
      p21_uge_8201 <= p21_data_enable ? p20_uge_8201 : p21_uge_8201;
      p21_uge_8283 <= p21_data_enable ? uge_8283 : p21_uge_8283;
      p21_concat_8288 <= p21_data_enable ? concat_8288 : p21_concat_8288;
      p21_uge_8289 <= p21_data_enable ? uge_8289 : p21_uge_8289;
      p21_bit_slice_6551 <= p21_data_enable ? p20_bit_slice_6551 : p21_bit_slice_6551;
      p21_bit_slice_6552 <= p21_data_enable ? p20_bit_slice_6552 : p21_bit_slice_6552;
      p21_bit_slice_6553 <= p21_data_enable ? p20_bit_slice_6553 : p21_bit_slice_6553;
      p21_bit_slice_6554 <= p21_data_enable ? p20_bit_slice_6554 : p21_bit_slice_6554;
      p21_bit_slice_6555 <= p21_data_enable ? p20_bit_slice_6555 : p21_bit_slice_6555;
      p21_negated <= p21_data_enable ? p20_negated : p21_negated;
      p22_b <= p22_data_enable ? p21_b : p22_b;
      p22_uge_6629 <= p22_data_enable ? p21_uge_6629 : p22_uge_6629;
      p22_bivisor__1 <= p22_data_enable ? p21_bivisor__1 : p22_bivisor__1;
      p22_uge_6637 <= p22_data_enable ? p21_uge_6637 : p22_uge_6637;
      p22_uge_6719 <= p22_data_enable ? p21_uge_6719 : p22_uge_6719;
      p22_uge_6801 <= p22_data_enable ? p21_uge_6801 : p22_uge_6801;
      p22_uge_6881 <= p22_data_enable ? p21_uge_6881 : p22_uge_6881;
      p22_uge_6963 <= p22_data_enable ? p21_uge_6963 : p22_uge_6963;
      p22_uge_6969 <= p22_data_enable ? p21_uge_6969 : p22_uge_6969;
      p22_uge_7049 <= p22_data_enable ? p21_uge_7049 : p22_uge_7049;
      p22_uge_7131 <= p22_data_enable ? p21_uge_7131 : p22_uge_7131;
      p22_uge_7211 <= p22_data_enable ? p21_uge_7211 : p22_uge_7211;
      p22_uge_7293 <= p22_data_enable ? p21_uge_7293 : p22_uge_7293;
      p22_uge_7299 <= p22_data_enable ? p21_uge_7299 : p22_uge_7299;
      p22_uge_7379 <= p22_data_enable ? p21_uge_7379 : p22_uge_7379;
      p22_uge_7461 <= p22_data_enable ? p21_uge_7461 : p22_uge_7461;
      p22_uge_7541 <= p22_data_enable ? p21_uge_7541 : p22_uge_7541;
      p22_uge_7623 <= p22_data_enable ? p21_uge_7623 : p22_uge_7623;
      p22_uge_7629 <= p22_data_enable ? p21_uge_7629 : p22_uge_7629;
      p22_uge_7709 <= p22_data_enable ? p21_uge_7709 : p22_uge_7709;
      p22_uge_7791 <= p22_data_enable ? p21_uge_7791 : p22_uge_7791;
      p22_uge_7871 <= p22_data_enable ? p21_uge_7871 : p22_uge_7871;
      p22_uge_7953 <= p22_data_enable ? p21_uge_7953 : p22_uge_7953;
      p22_uge_7959 <= p22_data_enable ? p21_uge_7959 : p22_uge_7959;
      p22_uge_8039 <= p22_data_enable ? p21_uge_8039 : p22_uge_8039;
      p22_uge_8121 <= p22_data_enable ? p21_uge_8121 : p22_uge_8121;
      p22_uge_8201 <= p22_data_enable ? p21_uge_8201 : p22_uge_8201;
      p22_uge_8283 <= p22_data_enable ? p21_uge_8283 : p22_uge_8283;
      p22_uge_8289 <= p22_data_enable ? p21_uge_8289 : p22_uge_8289;
      p22_concat_8368 <= p22_data_enable ? concat_8368 : p22_concat_8368;
      p22_uge_8369 <= p22_data_enable ? uge_8369 : p22_uge_8369;
      p22_sub_8370 <= p22_data_enable ? sub_8370 : p22_sub_8370;
      p22_bit_slice_6552 <= p22_data_enable ? p21_bit_slice_6552 : p22_bit_slice_6552;
      p22_bit_slice_6553 <= p22_data_enable ? p21_bit_slice_6553 : p22_bit_slice_6553;
      p22_bit_slice_6554 <= p22_data_enable ? p21_bit_slice_6554 : p22_bit_slice_6554;
      p22_bit_slice_6555 <= p22_data_enable ? p21_bit_slice_6555 : p22_bit_slice_6555;
      p22_negated <= p22_data_enable ? p21_negated : p22_negated;
      p23_b <= p23_data_enable ? p22_b : p23_b;
      p23_uge_6629 <= p23_data_enable ? p22_uge_6629 : p23_uge_6629;
      p23_bivisor__1 <= p23_data_enable ? p22_bivisor__1 : p23_bivisor__1;
      p23_uge_6637 <= p23_data_enable ? p22_uge_6637 : p23_uge_6637;
      p23_uge_6719 <= p23_data_enable ? p22_uge_6719 : p23_uge_6719;
      p23_uge_6801 <= p23_data_enable ? p22_uge_6801 : p23_uge_6801;
      p23_uge_6881 <= p23_data_enable ? p22_uge_6881 : p23_uge_6881;
      p23_uge_6963 <= p23_data_enable ? p22_uge_6963 : p23_uge_6963;
      p23_uge_6969 <= p23_data_enable ? p22_uge_6969 : p23_uge_6969;
      p23_uge_7049 <= p23_data_enable ? p22_uge_7049 : p23_uge_7049;
      p23_uge_7131 <= p23_data_enable ? p22_uge_7131 : p23_uge_7131;
      p23_uge_7211 <= p23_data_enable ? p22_uge_7211 : p23_uge_7211;
      p23_uge_7293 <= p23_data_enable ? p22_uge_7293 : p23_uge_7293;
      p23_uge_7299 <= p23_data_enable ? p22_uge_7299 : p23_uge_7299;
      p23_uge_7379 <= p23_data_enable ? p22_uge_7379 : p23_uge_7379;
      p23_uge_7461 <= p23_data_enable ? p22_uge_7461 : p23_uge_7461;
      p23_uge_7541 <= p23_data_enable ? p22_uge_7541 : p23_uge_7541;
      p23_uge_7623 <= p23_data_enable ? p22_uge_7623 : p23_uge_7623;
      p23_uge_7629 <= p23_data_enable ? p22_uge_7629 : p23_uge_7629;
      p23_uge_7709 <= p23_data_enable ? p22_uge_7709 : p23_uge_7709;
      p23_uge_7791 <= p23_data_enable ? p22_uge_7791 : p23_uge_7791;
      p23_uge_7871 <= p23_data_enable ? p22_uge_7871 : p23_uge_7871;
      p23_uge_7953 <= p23_data_enable ? p22_uge_7953 : p23_uge_7953;
      p23_uge_7959 <= p23_data_enable ? p22_uge_7959 : p23_uge_7959;
      p23_uge_8039 <= p23_data_enable ? p22_uge_8039 : p23_uge_8039;
      p23_uge_8121 <= p23_data_enable ? p22_uge_8121 : p23_uge_8121;
      p23_uge_8201 <= p23_data_enable ? p22_uge_8201 : p23_uge_8201;
      p23_uge_8283 <= p23_data_enable ? p22_uge_8283 : p23_uge_8283;
      p23_uge_8289 <= p23_data_enable ? p22_uge_8289 : p23_uge_8289;
      p23_uge_8369 <= p23_data_enable ? p22_uge_8369 : p23_uge_8369;
      p23_uge_8451 <= p23_data_enable ? uge_8451 : p23_uge_8451;
      p23_r__93 <= p23_data_enable ? r__93 : p23_r__93;
      p23_bit_slice_6553 <= p23_data_enable ? p22_bit_slice_6553 : p23_bit_slice_6553;
      p23_bit_slice_6554 <= p23_data_enable ? p22_bit_slice_6554 : p23_bit_slice_6554;
      p23_bit_slice_6555 <= p23_data_enable ? p22_bit_slice_6555 : p23_bit_slice_6555;
      p23_negated <= p23_data_enable ? p22_negated : p23_negated;
      p24_b <= p24_data_enable ? p23_b : p24_b;
      p24_uge_6629 <= p24_data_enable ? p23_uge_6629 : p24_uge_6629;
      p24_bivisor__1 <= p24_data_enable ? p23_bivisor__1 : p24_bivisor__1;
      p24_uge_6637 <= p24_data_enable ? p23_uge_6637 : p24_uge_6637;
      p24_uge_6719 <= p24_data_enable ? p23_uge_6719 : p24_uge_6719;
      p24_uge_6801 <= p24_data_enable ? p23_uge_6801 : p24_uge_6801;
      p24_uge_6881 <= p24_data_enable ? p23_uge_6881 : p24_uge_6881;
      p24_uge_6963 <= p24_data_enable ? p23_uge_6963 : p24_uge_6963;
      p24_uge_6969 <= p24_data_enable ? p23_uge_6969 : p24_uge_6969;
      p24_uge_7049 <= p24_data_enable ? p23_uge_7049 : p24_uge_7049;
      p24_uge_7131 <= p24_data_enable ? p23_uge_7131 : p24_uge_7131;
      p24_uge_7211 <= p24_data_enable ? p23_uge_7211 : p24_uge_7211;
      p24_uge_7293 <= p24_data_enable ? p23_uge_7293 : p24_uge_7293;
      p24_uge_7299 <= p24_data_enable ? p23_uge_7299 : p24_uge_7299;
      p24_uge_7379 <= p24_data_enable ? p23_uge_7379 : p24_uge_7379;
      p24_uge_7461 <= p24_data_enable ? p23_uge_7461 : p24_uge_7461;
      p24_uge_7541 <= p24_data_enable ? p23_uge_7541 : p24_uge_7541;
      p24_uge_7623 <= p24_data_enable ? p23_uge_7623 : p24_uge_7623;
      p24_uge_7629 <= p24_data_enable ? p23_uge_7629 : p24_uge_7629;
      p24_uge_7709 <= p24_data_enable ? p23_uge_7709 : p24_uge_7709;
      p24_uge_7791 <= p24_data_enable ? p23_uge_7791 : p24_uge_7791;
      p24_uge_7871 <= p24_data_enable ? p23_uge_7871 : p24_uge_7871;
      p24_uge_7953 <= p24_data_enable ? p23_uge_7953 : p24_uge_7953;
      p24_uge_7959 <= p24_data_enable ? p23_uge_7959 : p24_uge_7959;
      p24_uge_8039 <= p24_data_enable ? p23_uge_8039 : p24_uge_8039;
      p24_uge_8121 <= p24_data_enable ? p23_uge_8121 : p24_uge_8121;
      p24_uge_8201 <= p24_data_enable ? p23_uge_8201 : p24_uge_8201;
      p24_uge_8283 <= p24_data_enable ? p23_uge_8283 : p24_uge_8283;
      p24_uge_8289 <= p24_data_enable ? p23_uge_8289 : p24_uge_8289;
      p24_uge_8369 <= p24_data_enable ? p23_uge_8369 : p24_uge_8369;
      p24_uge_8451 <= p24_data_enable ? p23_uge_8451 : p24_uge_8451;
      p24_uge_8531 <= p24_data_enable ? uge_8531 : p24_uge_8531;
      p24_r__94 <= p24_data_enable ? r__94 : p24_r__94;
      p24_bit_slice_6554 <= p24_data_enable ? p23_bit_slice_6554 : p24_bit_slice_6554;
      p24_bit_slice_8534 <= p24_data_enable ? bit_slice_8534 : p24_bit_slice_8534;
      p24_bit_slice_6555 <= p24_data_enable ? p23_bit_slice_6555 : p24_bit_slice_6555;
      p24_negated <= p24_data_enable ? p23_negated : p24_negated;
      p25_uge_6629 <= p25_data_enable ? p24_uge_6629 : p25_uge_6629;
      p25_uge_6637 <= p25_data_enable ? p24_uge_6637 : p25_uge_6637;
      p25_uge_6719 <= p25_data_enable ? p24_uge_6719 : p25_uge_6719;
      p25_uge_6801 <= p25_data_enable ? p24_uge_6801 : p25_uge_6801;
      p25_uge_6881 <= p25_data_enable ? p24_uge_6881 : p25_uge_6881;
      p25_uge_6963 <= p25_data_enable ? p24_uge_6963 : p25_uge_6963;
      p25_uge_6969 <= p25_data_enable ? p24_uge_6969 : p25_uge_6969;
      p25_uge_7049 <= p25_data_enable ? p24_uge_7049 : p25_uge_7049;
      p25_uge_7131 <= p25_data_enable ? p24_uge_7131 : p25_uge_7131;
      p25_uge_7211 <= p25_data_enable ? p24_uge_7211 : p25_uge_7211;
      p25_uge_7293 <= p25_data_enable ? p24_uge_7293 : p25_uge_7293;
      p25_uge_7299 <= p25_data_enable ? p24_uge_7299 : p25_uge_7299;
      p25_uge_7379 <= p25_data_enable ? p24_uge_7379 : p25_uge_7379;
      p25_uge_7461 <= p25_data_enable ? p24_uge_7461 : p25_uge_7461;
      p25_uge_7541 <= p25_data_enable ? p24_uge_7541 : p25_uge_7541;
      p25_uge_7623 <= p25_data_enable ? p24_uge_7623 : p25_uge_7623;
      p25_uge_7629 <= p25_data_enable ? p24_uge_7629 : p25_uge_7629;
      p25_uge_7709 <= p25_data_enable ? p24_uge_7709 : p25_uge_7709;
      p25_uge_7791 <= p25_data_enable ? p24_uge_7791 : p25_uge_7791;
      p25_uge_7871 <= p25_data_enable ? p24_uge_7871 : p25_uge_7871;
      p25_uge_7953 <= p25_data_enable ? p24_uge_7953 : p25_uge_7953;
      p25_uge_7959 <= p25_data_enable ? p24_uge_7959 : p25_uge_7959;
      p25_uge_8039 <= p25_data_enable ? p24_uge_8039 : p25_uge_8039;
      p25_uge_8121 <= p25_data_enable ? p24_uge_8121 : p25_uge_8121;
      p25_uge_8201 <= p25_data_enable ? p24_uge_8201 : p25_uge_8201;
      p25_uge_8283 <= p25_data_enable ? p24_uge_8283 : p25_uge_8283;
      p25_uge_8289 <= p25_data_enable ? p24_uge_8289 : p25_uge_8289;
      p25_uge_8369 <= p25_data_enable ? p24_uge_8369 : p25_uge_8369;
      p25_uge_8451 <= p25_data_enable ? p24_uge_8451 : p25_uge_8451;
      p25_uge_8531 <= p25_data_enable ? p24_uge_8531 : p25_uge_8531;
      p25_uge_8613 <= p25_data_enable ? uge_8613 : p25_uge_8613;
      p25_q__32_squeezed_portion_0_width_1 <= p25_data_enable ? q__32_squeezed_portion_0_width_1 : p25_q__32_squeezed_portion_0_width_1;
      p25_negated <= p25_data_enable ? p24_negated : p25_negated;
      p0_valid <= p0_enable ? p0_all_active_inputs_valid : p0_valid;
      p1_valid <= p1_enable ? p0_valid : p1_valid;
      p2_valid <= p2_enable ? p1_valid : p2_valid;
      p3_valid <= p3_enable ? p2_valid : p3_valid;
      p4_valid <= p4_enable ? p3_valid : p4_valid;
      p5_valid <= p5_enable ? p4_valid : p5_valid;
      p6_valid <= p6_enable ? p5_valid : p6_valid;
      p7_valid <= p7_enable ? p6_valid : p7_valid;
      p8_valid <= p8_enable ? p7_valid : p8_valid;
      p9_valid <= p9_enable ? p8_valid : p9_valid;
      p10_valid <= p10_enable ? p9_valid : p10_valid;
      p11_valid <= p11_enable ? p10_valid : p11_valid;
      p12_valid <= p12_enable ? p11_valid : p12_valid;
      p13_valid <= p13_enable ? p12_valid : p13_valid;
      p14_valid <= p14_enable ? p13_valid : p14_valid;
      p15_valid <= p15_enable ? p14_valid : p15_valid;
      p16_valid <= p16_enable ? p15_valid : p16_valid;
      p17_valid <= p17_enable ? p16_valid : p17_valid;
      p18_valid <= p18_enable ? p17_valid : p18_valid;
      p19_valid <= p19_enable ? p18_valid : p19_valid;
      p20_valid <= p20_enable ? p19_valid : p20_valid;
      p21_valid <= p21_enable ? p20_valid : p21_valid;
      p22_valid <= p22_enable ? p21_valid : p22_valid;
      p23_valid <= p23_enable ? p22_valid : p23_valid;
      p24_valid <= p24_enable ? p23_valid : p24_valid;
      p25_valid <= p25_enable ? p24_valid : p25_valid;
      p26_valid <= p26_enable ? p26_stage_done : p26_valid;
      p27_valid <= p27_enable ? p26_valid : p27_valid;
      p28_valid <= p28_enable ? p27_valid : p28_valid;
      p29_valid <= p29_enable ? p28_valid : p29_valid;
      p30_valid <= p30_enable ? p29_valid : p30_valid;
      lhs_reg <= lhs_load_en ? lhs : lhs_reg;
      lhs_valid_reg <= lhs_valid_load_en ? lhs_valid : lhs_valid_reg;
      rhs_reg <= rhs_load_en ? rhs : rhs_reg;
      rhs_valid_reg <= rhs_valid_load_en ? rhs_valid : rhs_valid_reg;
      result_reg <= result_load_en ? signed_div : result_reg;
      result_valid_reg <= result_valid_load_en ? p25_valid : result_valid_reg;
    end
  end
  assign result = result_reg;
  assign result_valid = result_valid_reg;
  assign lhs_ready = lhs_load_en;
  assign rhs_ready = rhs_load_en;
endmodule
module xls_divui32(
  input wire clk,
  input wire rst,
  input wire [31:0] lhs,
  input wire lhs_valid,
  input wire [31:0] rhs,
  input wire rhs_valid,
  input wire result_ready,
  output wire [31:0] result,
  output wire result_valid,
  output wire lhs_ready,
  output wire rhs_ready
);
  reg [31:0] p0_concat_6500;
  reg [31:0] p0_b;
  reg p0_uge_6502;
  reg [31:0] p0_sub_6503;
  reg p0_bit_slice_6504;
  reg p0_bit_slice_6505;
  reg p0_bit_slice_6506;
  reg p0_bit_slice_6507;
  reg p0_bit_slice_6508;
  reg p0_bit_slice_6509;
  reg p0_bit_slice_6510;
  reg p0_bit_slice_6511;
  reg p0_bit_slice_6512;
  reg p0_bit_slice_6513;
  reg p0_bit_slice_6514;
  reg p0_bit_slice_6515;
  reg p0_bit_slice_6516;
  reg p0_bit_slice_6517;
  reg p0_bit_slice_6518;
  reg p0_bit_slice_6519;
  reg p0_bit_slice_6520;
  reg p0_bit_slice_6521;
  reg p0_bit_slice_6522;
  reg p0_bit_slice_6523;
  reg p0_bit_slice_6524;
  reg p0_bit_slice_6525;
  reg p0_bit_slice_6526;
  reg p0_bit_slice_6527;
  reg p0_bit_slice_6528;
  reg p0_bit_slice_6529;
  reg p0_bit_slice_6530;
  reg p0_bit_slice_6531;
  reg p0_bit_slice_6532;
  reg p0_bit_slice_6533;
  reg p0_bit_slice_6534;
  reg [31:0] p1_b;
  reg p1_uge_6502;
  reg [32:0] p1_bivisor__1;
  reg p1_uge_6616;
  reg [31:0] p1_r__66;
  reg p1_bit_slice_6505;
  reg p1_bit_slice_6506;
  reg p1_bit_slice_6507;
  reg p1_bit_slice_6508;
  reg p1_bit_slice_6509;
  reg p1_bit_slice_6510;
  reg p1_bit_slice_6511;
  reg p1_bit_slice_6512;
  reg p1_bit_slice_6513;
  reg p1_bit_slice_6514;
  reg p1_bit_slice_6515;
  reg p1_bit_slice_6516;
  reg p1_bit_slice_6517;
  reg p1_bit_slice_6518;
  reg p1_bit_slice_6519;
  reg p1_bit_slice_6520;
  reg p1_bit_slice_6521;
  reg p1_bit_slice_6522;
  reg p1_bit_slice_6523;
  reg p1_bit_slice_6524;
  reg p1_bit_slice_6525;
  reg p1_bit_slice_6526;
  reg p1_bit_slice_6527;
  reg p1_bit_slice_6528;
  reg p1_bit_slice_6529;
  reg p1_bit_slice_6530;
  reg p1_bit_slice_6531;
  reg p1_bit_slice_6532;
  reg p1_bit_slice_6533;
  reg p1_bit_slice_6534;
  reg [31:0] p2_b;
  reg p2_uge_6502;
  reg [32:0] p2_bivisor__1;
  reg p2_uge_6616;
  reg p2_uge_6694;
  reg [31:0] p2_r__67;
  reg p2_bit_slice_6506;
  reg [30:0] p2_bit_slice_6697;
  reg p2_bit_slice_6507;
  reg p2_bit_slice_6508;
  reg p2_bit_slice_6509;
  reg p2_bit_slice_6510;
  reg p2_bit_slice_6511;
  reg p2_bit_slice_6512;
  reg p2_bit_slice_6513;
  reg p2_bit_slice_6514;
  reg p2_bit_slice_6515;
  reg p2_bit_slice_6516;
  reg p2_bit_slice_6517;
  reg p2_bit_slice_6518;
  reg p2_bit_slice_6519;
  reg p2_bit_slice_6520;
  reg p2_bit_slice_6521;
  reg p2_bit_slice_6522;
  reg p2_bit_slice_6523;
  reg p2_bit_slice_6524;
  reg p2_bit_slice_6525;
  reg p2_bit_slice_6526;
  reg p2_bit_slice_6527;
  reg p2_bit_slice_6528;
  reg p2_bit_slice_6529;
  reg p2_bit_slice_6530;
  reg p2_bit_slice_6531;
  reg p2_bit_slice_6532;
  reg p2_bit_slice_6533;
  reg p2_bit_slice_6534;
  reg [31:0] p3_b;
  reg p3_uge_6502;
  reg [32:0] p3_bivisor__1;
  reg p3_uge_6616;
  reg p3_uge_6694;
  reg p3_uge_6774;
  reg [31:0] p3_concat_6779;
  reg p3_uge_6780;
  reg p3_bit_slice_6508;
  reg p3_bit_slice_6509;
  reg p3_bit_slice_6510;
  reg p3_bit_slice_6511;
  reg p3_bit_slice_6512;
  reg p3_bit_slice_6513;
  reg p3_bit_slice_6514;
  reg p3_bit_slice_6515;
  reg p3_bit_slice_6516;
  reg p3_bit_slice_6517;
  reg p3_bit_slice_6518;
  reg p3_bit_slice_6519;
  reg p3_bit_slice_6520;
  reg p3_bit_slice_6521;
  reg p3_bit_slice_6522;
  reg p3_bit_slice_6523;
  reg p3_bit_slice_6524;
  reg p3_bit_slice_6525;
  reg p3_bit_slice_6526;
  reg p3_bit_slice_6527;
  reg p3_bit_slice_6528;
  reg p3_bit_slice_6529;
  reg p3_bit_slice_6530;
  reg p3_bit_slice_6531;
  reg p3_bit_slice_6532;
  reg p3_bit_slice_6533;
  reg p3_bit_slice_6534;
  reg [31:0] p4_b;
  reg p4_uge_6502;
  reg [32:0] p4_bivisor__1;
  reg p4_uge_6616;
  reg p4_uge_6694;
  reg p4_uge_6774;
  reg p4_uge_6780;
  reg [31:0] p4_concat_6857;
  reg p4_uge_6858;
  reg [31:0] p4_sub_6859;
  reg p4_bit_slice_6509;
  reg p4_bit_slice_6510;
  reg p4_bit_slice_6511;
  reg p4_bit_slice_6512;
  reg p4_bit_slice_6513;
  reg p4_bit_slice_6514;
  reg p4_bit_slice_6515;
  reg p4_bit_slice_6516;
  reg p4_bit_slice_6517;
  reg p4_bit_slice_6518;
  reg p4_bit_slice_6519;
  reg p4_bit_slice_6520;
  reg p4_bit_slice_6521;
  reg p4_bit_slice_6522;
  reg p4_bit_slice_6523;
  reg p4_bit_slice_6524;
  reg p4_bit_slice_6525;
  reg p4_bit_slice_6526;
  reg p4_bit_slice_6527;
  reg p4_bit_slice_6528;
  reg p4_bit_slice_6529;
  reg p4_bit_slice_6530;
  reg p4_bit_slice_6531;
  reg p4_bit_slice_6532;
  reg p4_bit_slice_6533;
  reg p4_bit_slice_6534;
  reg [31:0] p5_b;
  reg p5_uge_6502;
  reg [32:0] p5_bivisor__1;
  reg p5_uge_6616;
  reg p5_uge_6694;
  reg p5_uge_6774;
  reg p5_uge_6780;
  reg p5_uge_6858;
  reg p5_uge_6938;
  reg [31:0] p5_r__71;
  reg p5_bit_slice_6510;
  reg p5_bit_slice_6511;
  reg p5_bit_slice_6512;
  reg p5_bit_slice_6513;
  reg p5_bit_slice_6514;
  reg p5_bit_slice_6515;
  reg p5_bit_slice_6516;
  reg p5_bit_slice_6517;
  reg p5_bit_slice_6518;
  reg p5_bit_slice_6519;
  reg p5_bit_slice_6520;
  reg p5_bit_slice_6521;
  reg p5_bit_slice_6522;
  reg p5_bit_slice_6523;
  reg p5_bit_slice_6524;
  reg p5_bit_slice_6525;
  reg p5_bit_slice_6526;
  reg p5_bit_slice_6527;
  reg p5_bit_slice_6528;
  reg p5_bit_slice_6529;
  reg p5_bit_slice_6530;
  reg p5_bit_slice_6531;
  reg p5_bit_slice_6532;
  reg p5_bit_slice_6533;
  reg p5_bit_slice_6534;
  reg [31:0] p6_b;
  reg p6_uge_6502;
  reg [32:0] p6_bivisor__1;
  reg p6_uge_6616;
  reg p6_uge_6694;
  reg p6_uge_6774;
  reg p6_uge_6780;
  reg p6_uge_6858;
  reg p6_uge_6938;
  reg p6_uge_7016;
  reg [31:0] p6_r__72;
  reg p6_bit_slice_6511;
  reg [30:0] p6_bit_slice_7019;
  reg p6_bit_slice_6512;
  reg p6_bit_slice_6513;
  reg p6_bit_slice_6514;
  reg p6_bit_slice_6515;
  reg p6_bit_slice_6516;
  reg p6_bit_slice_6517;
  reg p6_bit_slice_6518;
  reg p6_bit_slice_6519;
  reg p6_bit_slice_6520;
  reg p6_bit_slice_6521;
  reg p6_bit_slice_6522;
  reg p6_bit_slice_6523;
  reg p6_bit_slice_6524;
  reg p6_bit_slice_6525;
  reg p6_bit_slice_6526;
  reg p6_bit_slice_6527;
  reg p6_bit_slice_6528;
  reg p6_bit_slice_6529;
  reg p6_bit_slice_6530;
  reg p6_bit_slice_6531;
  reg p6_bit_slice_6532;
  reg p6_bit_slice_6533;
  reg p6_bit_slice_6534;
  reg [31:0] p7_b;
  reg p7_uge_6502;
  reg [32:0] p7_bivisor__1;
  reg p7_uge_6616;
  reg p7_uge_6694;
  reg p7_uge_6774;
  reg p7_uge_6780;
  reg p7_uge_6858;
  reg p7_uge_6938;
  reg p7_uge_7016;
  reg p7_uge_7096;
  reg [31:0] p7_concat_7101;
  reg p7_uge_7102;
  reg p7_bit_slice_6513;
  reg p7_bit_slice_6514;
  reg p7_bit_slice_6515;
  reg p7_bit_slice_6516;
  reg p7_bit_slice_6517;
  reg p7_bit_slice_6518;
  reg p7_bit_slice_6519;
  reg p7_bit_slice_6520;
  reg p7_bit_slice_6521;
  reg p7_bit_slice_6522;
  reg p7_bit_slice_6523;
  reg p7_bit_slice_6524;
  reg p7_bit_slice_6525;
  reg p7_bit_slice_6526;
  reg p7_bit_slice_6527;
  reg p7_bit_slice_6528;
  reg p7_bit_slice_6529;
  reg p7_bit_slice_6530;
  reg p7_bit_slice_6531;
  reg p7_bit_slice_6532;
  reg p7_bit_slice_6533;
  reg p7_bit_slice_6534;
  reg [31:0] p8_b;
  reg p8_uge_6502;
  reg [32:0] p8_bivisor__1;
  reg p8_uge_6616;
  reg p8_uge_6694;
  reg p8_uge_6774;
  reg p8_uge_6780;
  reg p8_uge_6858;
  reg p8_uge_6938;
  reg p8_uge_7016;
  reg p8_uge_7096;
  reg p8_uge_7102;
  reg [31:0] p8_concat_7179;
  reg p8_uge_7180;
  reg [31:0] p8_sub_7181;
  reg p8_bit_slice_6514;
  reg p8_bit_slice_6515;
  reg p8_bit_slice_6516;
  reg p8_bit_slice_6517;
  reg p8_bit_slice_6518;
  reg p8_bit_slice_6519;
  reg p8_bit_slice_6520;
  reg p8_bit_slice_6521;
  reg p8_bit_slice_6522;
  reg p8_bit_slice_6523;
  reg p8_bit_slice_6524;
  reg p8_bit_slice_6525;
  reg p8_bit_slice_6526;
  reg p8_bit_slice_6527;
  reg p8_bit_slice_6528;
  reg p8_bit_slice_6529;
  reg p8_bit_slice_6530;
  reg p8_bit_slice_6531;
  reg p8_bit_slice_6532;
  reg p8_bit_slice_6533;
  reg p8_bit_slice_6534;
  reg [31:0] p9_b;
  reg p9_uge_6502;
  reg [32:0] p9_bivisor__1;
  reg p9_uge_6616;
  reg p9_uge_6694;
  reg p9_uge_6774;
  reg p9_uge_6780;
  reg p9_uge_6858;
  reg p9_uge_6938;
  reg p9_uge_7016;
  reg p9_uge_7096;
  reg p9_uge_7102;
  reg p9_uge_7180;
  reg p9_uge_7260;
  reg [31:0] p9_r__76;
  reg p9_bit_slice_6515;
  reg p9_bit_slice_6516;
  reg p9_bit_slice_6517;
  reg p9_bit_slice_6518;
  reg p9_bit_slice_6519;
  reg p9_bit_slice_6520;
  reg p9_bit_slice_6521;
  reg p9_bit_slice_6522;
  reg p9_bit_slice_6523;
  reg p9_bit_slice_6524;
  reg p9_bit_slice_6525;
  reg p9_bit_slice_6526;
  reg p9_bit_slice_6527;
  reg p9_bit_slice_6528;
  reg p9_bit_slice_6529;
  reg p9_bit_slice_6530;
  reg p9_bit_slice_6531;
  reg p9_bit_slice_6532;
  reg p9_bit_slice_6533;
  reg p9_bit_slice_6534;
  reg [31:0] p10_b;
  reg p10_uge_6502;
  reg [32:0] p10_bivisor__1;
  reg p10_uge_6616;
  reg p10_uge_6694;
  reg p10_uge_6774;
  reg p10_uge_6780;
  reg p10_uge_6858;
  reg p10_uge_6938;
  reg p10_uge_7016;
  reg p10_uge_7096;
  reg p10_uge_7102;
  reg p10_uge_7180;
  reg p10_uge_7260;
  reg p10_uge_7338;
  reg [31:0] p10_r__77;
  reg p10_bit_slice_6516;
  reg [30:0] p10_bit_slice_7341;
  reg p10_bit_slice_6517;
  reg p10_bit_slice_6518;
  reg p10_bit_slice_6519;
  reg p10_bit_slice_6520;
  reg p10_bit_slice_6521;
  reg p10_bit_slice_6522;
  reg p10_bit_slice_6523;
  reg p10_bit_slice_6524;
  reg p10_bit_slice_6525;
  reg p10_bit_slice_6526;
  reg p10_bit_slice_6527;
  reg p10_bit_slice_6528;
  reg p10_bit_slice_6529;
  reg p10_bit_slice_6530;
  reg p10_bit_slice_6531;
  reg p10_bit_slice_6532;
  reg p10_bit_slice_6533;
  reg p10_bit_slice_6534;
  reg [31:0] p11_b;
  reg p11_uge_6502;
  reg [32:0] p11_bivisor__1;
  reg p11_uge_6616;
  reg p11_uge_6694;
  reg p11_uge_6774;
  reg p11_uge_6780;
  reg p11_uge_6858;
  reg p11_uge_6938;
  reg p11_uge_7016;
  reg p11_uge_7096;
  reg p11_uge_7102;
  reg p11_uge_7180;
  reg p11_uge_7260;
  reg p11_uge_7338;
  reg p11_uge_7418;
  reg [31:0] p11_concat_7423;
  reg p11_uge_7424;
  reg p11_bit_slice_6518;
  reg p11_bit_slice_6519;
  reg p11_bit_slice_6520;
  reg p11_bit_slice_6521;
  reg p11_bit_slice_6522;
  reg p11_bit_slice_6523;
  reg p11_bit_slice_6524;
  reg p11_bit_slice_6525;
  reg p11_bit_slice_6526;
  reg p11_bit_slice_6527;
  reg p11_bit_slice_6528;
  reg p11_bit_slice_6529;
  reg p11_bit_slice_6530;
  reg p11_bit_slice_6531;
  reg p11_bit_slice_6532;
  reg p11_bit_slice_6533;
  reg p11_bit_slice_6534;
  reg [31:0] p12_b;
  reg p12_uge_6502;
  reg [32:0] p12_bivisor__1;
  reg p12_uge_6616;
  reg p12_uge_6694;
  reg p12_uge_6774;
  reg p12_uge_6780;
  reg p12_uge_6858;
  reg p12_uge_6938;
  reg p12_uge_7016;
  reg p12_uge_7096;
  reg p12_uge_7102;
  reg p12_uge_7180;
  reg p12_uge_7260;
  reg p12_uge_7338;
  reg p12_uge_7418;
  reg p12_uge_7424;
  reg [31:0] p12_concat_7501;
  reg p12_uge_7502;
  reg [31:0] p12_sub_7503;
  reg p12_bit_slice_6519;
  reg p12_bit_slice_6520;
  reg p12_bit_slice_6521;
  reg p12_bit_slice_6522;
  reg p12_bit_slice_6523;
  reg p12_bit_slice_6524;
  reg p12_bit_slice_6525;
  reg p12_bit_slice_6526;
  reg p12_bit_slice_6527;
  reg p12_bit_slice_6528;
  reg p12_bit_slice_6529;
  reg p12_bit_slice_6530;
  reg p12_bit_slice_6531;
  reg p12_bit_slice_6532;
  reg p12_bit_slice_6533;
  reg p12_bit_slice_6534;
  reg [31:0] p13_b;
  reg p13_uge_6502;
  reg [32:0] p13_bivisor__1;
  reg p13_uge_6616;
  reg p13_uge_6694;
  reg p13_uge_6774;
  reg p13_uge_6780;
  reg p13_uge_6858;
  reg p13_uge_6938;
  reg p13_uge_7016;
  reg p13_uge_7096;
  reg p13_uge_7102;
  reg p13_uge_7180;
  reg p13_uge_7260;
  reg p13_uge_7338;
  reg p13_uge_7418;
  reg p13_uge_7424;
  reg p13_uge_7502;
  reg p13_uge_7582;
  reg [31:0] p13_r__81;
  reg p13_bit_slice_6520;
  reg p13_bit_slice_6521;
  reg p13_bit_slice_6522;
  reg p13_bit_slice_6523;
  reg p13_bit_slice_6524;
  reg p13_bit_slice_6525;
  reg p13_bit_slice_6526;
  reg p13_bit_slice_6527;
  reg p13_bit_slice_6528;
  reg p13_bit_slice_6529;
  reg p13_bit_slice_6530;
  reg p13_bit_slice_6531;
  reg p13_bit_slice_6532;
  reg p13_bit_slice_6533;
  reg p13_bit_slice_6534;
  reg [31:0] p14_b;
  reg p14_uge_6502;
  reg [32:0] p14_bivisor__1;
  reg p14_uge_6616;
  reg p14_uge_6694;
  reg p14_uge_6774;
  reg p14_uge_6780;
  reg p14_uge_6858;
  reg p14_uge_6938;
  reg p14_uge_7016;
  reg p14_uge_7096;
  reg p14_uge_7102;
  reg p14_uge_7180;
  reg p14_uge_7260;
  reg p14_uge_7338;
  reg p14_uge_7418;
  reg p14_uge_7424;
  reg p14_uge_7502;
  reg p14_uge_7582;
  reg p14_uge_7660;
  reg [31:0] p14_r__82;
  reg p14_bit_slice_6521;
  reg [30:0] p14_bit_slice_7663;
  reg p14_bit_slice_6522;
  reg p14_bit_slice_6523;
  reg p14_bit_slice_6524;
  reg p14_bit_slice_6525;
  reg p14_bit_slice_6526;
  reg p14_bit_slice_6527;
  reg p14_bit_slice_6528;
  reg p14_bit_slice_6529;
  reg p14_bit_slice_6530;
  reg p14_bit_slice_6531;
  reg p14_bit_slice_6532;
  reg p14_bit_slice_6533;
  reg p14_bit_slice_6534;
  reg [31:0] p15_b;
  reg p15_uge_6502;
  reg [32:0] p15_bivisor__1;
  reg p15_uge_6616;
  reg p15_uge_6694;
  reg p15_uge_6774;
  reg p15_uge_6780;
  reg p15_uge_6858;
  reg p15_uge_6938;
  reg p15_uge_7016;
  reg p15_uge_7096;
  reg p15_uge_7102;
  reg p15_uge_7180;
  reg p15_uge_7260;
  reg p15_uge_7338;
  reg p15_uge_7418;
  reg p15_uge_7424;
  reg p15_uge_7502;
  reg p15_uge_7582;
  reg p15_uge_7660;
  reg p15_uge_7740;
  reg [31:0] p15_concat_7745;
  reg p15_uge_7746;
  reg p15_bit_slice_6523;
  reg p15_bit_slice_6524;
  reg p15_bit_slice_6525;
  reg p15_bit_slice_6526;
  reg p15_bit_slice_6527;
  reg p15_bit_slice_6528;
  reg p15_bit_slice_6529;
  reg p15_bit_slice_6530;
  reg p15_bit_slice_6531;
  reg p15_bit_slice_6532;
  reg p15_bit_slice_6533;
  reg p15_bit_slice_6534;
  reg [31:0] p16_b;
  reg p16_uge_6502;
  reg [32:0] p16_bivisor__1;
  reg p16_uge_6616;
  reg p16_uge_6694;
  reg p16_uge_6774;
  reg p16_uge_6780;
  reg p16_uge_6858;
  reg p16_uge_6938;
  reg p16_uge_7016;
  reg p16_uge_7096;
  reg p16_uge_7102;
  reg p16_uge_7180;
  reg p16_uge_7260;
  reg p16_uge_7338;
  reg p16_uge_7418;
  reg p16_uge_7424;
  reg p16_uge_7502;
  reg p16_uge_7582;
  reg p16_uge_7660;
  reg p16_uge_7740;
  reg p16_uge_7746;
  reg [31:0] p16_concat_7823;
  reg p16_uge_7824;
  reg [31:0] p16_sub_7825;
  reg p16_bit_slice_6524;
  reg p16_bit_slice_6525;
  reg p16_bit_slice_6526;
  reg p16_bit_slice_6527;
  reg p16_bit_slice_6528;
  reg p16_bit_slice_6529;
  reg p16_bit_slice_6530;
  reg p16_bit_slice_6531;
  reg p16_bit_slice_6532;
  reg p16_bit_slice_6533;
  reg p16_bit_slice_6534;
  reg [31:0] p17_b;
  reg p17_uge_6502;
  reg [32:0] p17_bivisor__1;
  reg p17_uge_6616;
  reg p17_uge_6694;
  reg p17_uge_6774;
  reg p17_uge_6780;
  reg p17_uge_6858;
  reg p17_uge_6938;
  reg p17_uge_7016;
  reg p17_uge_7096;
  reg p17_uge_7102;
  reg p17_uge_7180;
  reg p17_uge_7260;
  reg p17_uge_7338;
  reg p17_uge_7418;
  reg p17_uge_7424;
  reg p17_uge_7502;
  reg p17_uge_7582;
  reg p17_uge_7660;
  reg p17_uge_7740;
  reg p17_uge_7746;
  reg p17_uge_7824;
  reg p17_uge_7904;
  reg [31:0] p17_r__86;
  reg p17_bit_slice_6525;
  reg p17_bit_slice_6526;
  reg p17_bit_slice_6527;
  reg p17_bit_slice_6528;
  reg p17_bit_slice_6529;
  reg p17_bit_slice_6530;
  reg p17_bit_slice_6531;
  reg p17_bit_slice_6532;
  reg p17_bit_slice_6533;
  reg p17_bit_slice_6534;
  reg [31:0] p18_b;
  reg p18_uge_6502;
  reg [32:0] p18_bivisor__1;
  reg p18_uge_6616;
  reg p18_uge_6694;
  reg p18_uge_6774;
  reg p18_uge_6780;
  reg p18_uge_6858;
  reg p18_uge_6938;
  reg p18_uge_7016;
  reg p18_uge_7096;
  reg p18_uge_7102;
  reg p18_uge_7180;
  reg p18_uge_7260;
  reg p18_uge_7338;
  reg p18_uge_7418;
  reg p18_uge_7424;
  reg p18_uge_7502;
  reg p18_uge_7582;
  reg p18_uge_7660;
  reg p18_uge_7740;
  reg p18_uge_7746;
  reg p18_uge_7824;
  reg p18_uge_7904;
  reg p18_uge_7982;
  reg [31:0] p18_r__87;
  reg p18_bit_slice_6526;
  reg [30:0] p18_bit_slice_7985;
  reg p18_bit_slice_6527;
  reg p18_bit_slice_6528;
  reg p18_bit_slice_6529;
  reg p18_bit_slice_6530;
  reg p18_bit_slice_6531;
  reg p18_bit_slice_6532;
  reg p18_bit_slice_6533;
  reg p18_bit_slice_6534;
  reg [31:0] p19_b;
  reg p19_uge_6502;
  reg [32:0] p19_bivisor__1;
  reg p19_uge_6616;
  reg p19_uge_6694;
  reg p19_uge_6774;
  reg p19_uge_6780;
  reg p19_uge_6858;
  reg p19_uge_6938;
  reg p19_uge_7016;
  reg p19_uge_7096;
  reg p19_uge_7102;
  reg p19_uge_7180;
  reg p19_uge_7260;
  reg p19_uge_7338;
  reg p19_uge_7418;
  reg p19_uge_7424;
  reg p19_uge_7502;
  reg p19_uge_7582;
  reg p19_uge_7660;
  reg p19_uge_7740;
  reg p19_uge_7746;
  reg p19_uge_7824;
  reg p19_uge_7904;
  reg p19_uge_7982;
  reg p19_uge_8062;
  reg [31:0] p19_concat_8067;
  reg p19_uge_8068;
  reg p19_bit_slice_6528;
  reg p19_bit_slice_6529;
  reg p19_bit_slice_6530;
  reg p19_bit_slice_6531;
  reg p19_bit_slice_6532;
  reg p19_bit_slice_6533;
  reg p19_bit_slice_6534;
  reg [31:0] p20_b;
  reg p20_uge_6502;
  reg [32:0] p20_bivisor__1;
  reg p20_uge_6616;
  reg p20_uge_6694;
  reg p20_uge_6774;
  reg p20_uge_6780;
  reg p20_uge_6858;
  reg p20_uge_6938;
  reg p20_uge_7016;
  reg p20_uge_7096;
  reg p20_uge_7102;
  reg p20_uge_7180;
  reg p20_uge_7260;
  reg p20_uge_7338;
  reg p20_uge_7418;
  reg p20_uge_7424;
  reg p20_uge_7502;
  reg p20_uge_7582;
  reg p20_uge_7660;
  reg p20_uge_7740;
  reg p20_uge_7746;
  reg p20_uge_7824;
  reg p20_uge_7904;
  reg p20_uge_7982;
  reg p20_uge_8062;
  reg p20_uge_8068;
  reg [31:0] p20_concat_8145;
  reg p20_uge_8146;
  reg [31:0] p20_sub_8147;
  reg p20_bit_slice_6529;
  reg p20_bit_slice_6530;
  reg p20_bit_slice_6531;
  reg p20_bit_slice_6532;
  reg p20_bit_slice_6533;
  reg p20_bit_slice_6534;
  reg [31:0] p21_b;
  reg p21_uge_6502;
  reg [32:0] p21_bivisor__1;
  reg p21_uge_6616;
  reg p21_uge_6694;
  reg p21_uge_6774;
  reg p21_uge_6780;
  reg p21_uge_6858;
  reg p21_uge_6938;
  reg p21_uge_7016;
  reg p21_uge_7096;
  reg p21_uge_7102;
  reg p21_uge_7180;
  reg p21_uge_7260;
  reg p21_uge_7338;
  reg p21_uge_7418;
  reg p21_uge_7424;
  reg p21_uge_7502;
  reg p21_uge_7582;
  reg p21_uge_7660;
  reg p21_uge_7740;
  reg p21_uge_7746;
  reg p21_uge_7824;
  reg p21_uge_7904;
  reg p21_uge_7982;
  reg p21_uge_8062;
  reg p21_uge_8068;
  reg p21_uge_8146;
  reg p21_uge_8226;
  reg [31:0] p21_r__91;
  reg p21_bit_slice_6530;
  reg p21_bit_slice_6531;
  reg p21_bit_slice_6532;
  reg p21_bit_slice_6533;
  reg p21_bit_slice_6534;
  reg [31:0] p22_b;
  reg p22_uge_6502;
  reg [32:0] p22_bivisor__1;
  reg p22_uge_6616;
  reg p22_uge_6694;
  reg p22_uge_6774;
  reg p22_uge_6780;
  reg p22_uge_6858;
  reg p22_uge_6938;
  reg p22_uge_7016;
  reg p22_uge_7096;
  reg p22_uge_7102;
  reg p22_uge_7180;
  reg p22_uge_7260;
  reg p22_uge_7338;
  reg p22_uge_7418;
  reg p22_uge_7424;
  reg p22_uge_7502;
  reg p22_uge_7582;
  reg p22_uge_7660;
  reg p22_uge_7740;
  reg p22_uge_7746;
  reg p22_uge_7824;
  reg p22_uge_7904;
  reg p22_uge_7982;
  reg p22_uge_8062;
  reg p22_uge_8068;
  reg p22_uge_8146;
  reg p22_uge_8226;
  reg p22_uge_8304;
  reg [31:0] p22_r__92;
  reg p22_bit_slice_6531;
  reg [30:0] p22_bit_slice_8307;
  reg p22_bit_slice_6532;
  reg p22_bit_slice_6533;
  reg p22_bit_slice_6534;
  reg [31:0] p23_b;
  reg p23_uge_6502;
  reg [32:0] p23_bivisor__1;
  reg p23_uge_6616;
  reg p23_uge_6694;
  reg p23_uge_6774;
  reg p23_uge_6780;
  reg p23_uge_6858;
  reg p23_uge_6938;
  reg p23_uge_7016;
  reg p23_uge_7096;
  reg p23_uge_7102;
  reg p23_uge_7180;
  reg p23_uge_7260;
  reg p23_uge_7338;
  reg p23_uge_7418;
  reg p23_uge_7424;
  reg p23_uge_7502;
  reg p23_uge_7582;
  reg p23_uge_7660;
  reg p23_uge_7740;
  reg p23_uge_7746;
  reg p23_uge_7824;
  reg p23_uge_7904;
  reg p23_uge_7982;
  reg p23_uge_8062;
  reg p23_uge_8068;
  reg p23_uge_8146;
  reg p23_uge_8226;
  reg p23_uge_8304;
  reg p23_uge_8384;
  reg [31:0] p23_concat_8389;
  reg p23_uge_8390;
  reg p23_bit_slice_6533;
  reg p23_bit_slice_6534;
  reg p24_uge_6502;
  reg [32:0] p24_bivisor__1;
  reg p24_uge_6616;
  reg p24_uge_6694;
  reg p24_uge_6774;
  reg p24_uge_6780;
  reg p24_uge_6858;
  reg p24_uge_6938;
  reg p24_uge_7016;
  reg p24_uge_7096;
  reg p24_uge_7102;
  reg p24_uge_7180;
  reg p24_uge_7260;
  reg p24_uge_7338;
  reg p24_uge_7418;
  reg p24_uge_7424;
  reg p24_uge_7502;
  reg p24_uge_7582;
  reg p24_uge_7660;
  reg p24_uge_7740;
  reg p24_uge_7746;
  reg p24_uge_7824;
  reg p24_uge_7904;
  reg p24_uge_7982;
  reg p24_uge_8062;
  reg p24_uge_8068;
  reg p24_uge_8146;
  reg p24_uge_8226;
  reg p24_uge_8304;
  reg p24_uge_8384;
  reg p24_uge_8390;
  reg [31:0] p24_concat_8467;
  reg p24_uge_8468;
  reg [31:0] p24_sub_8469;
  reg p24_bit_slice_6534;
  reg p0_valid;
  reg p1_valid;
  reg p2_valid;
  reg p3_valid;
  reg p4_valid;
  reg p5_valid;
  reg p6_valid;
  reg p7_valid;
  reg p8_valid;
  reg p9_valid;
  reg p10_valid;
  reg p11_valid;
  reg p12_valid;
  reg p13_valid;
  reg p14_valid;
  reg p15_valid;
  reg p16_valid;
  reg p17_valid;
  reg p18_valid;
  reg p19_valid;
  reg p20_valid;
  reg p21_valid;
  reg p22_valid;
  reg p23_valid;
  reg p24_valid;
  reg p25_valid;
  reg p26_valid;
  reg p27_valid;
  reg p28_valid;
  reg p29_valid;
  reg p30_valid;
  reg [31:0] lhs_reg;
  reg lhs_valid_reg;
  reg [31:0] rhs_reg;
  reg rhs_valid_reg;
  reg [31:0] result_reg;
  reg result_valid_reg;
  wire result_valid_inv;
  wire result_valid_load_en;
  wire result_load_en;
  wire p25_stage_done;
  wire p25_not_valid;
  wire p24_enable;
  wire p24_data_enable;
  wire p24_not_valid;
  wire p23_enable;
  wire p23_data_enable;
  wire p23_not_valid;
  wire p22_enable;
  wire p22_data_enable;
  wire p22_not_valid;
  wire p21_enable;
  wire p21_data_enable;
  wire p21_not_valid;
  wire p20_enable;
  wire p20_data_enable;
  wire p20_not_valid;
  wire p19_enable;
  wire p19_data_enable;
  wire p19_not_valid;
  wire p18_enable;
  wire p18_data_enable;
  wire p18_not_valid;
  wire p17_enable;
  wire p17_data_enable;
  wire p17_not_valid;
  wire p16_enable;
  wire p16_data_enable;
  wire p16_not_valid;
  wire p15_enable;
  wire p15_data_enable;
  wire p15_not_valid;
  wire p14_enable;
  wire p14_data_enable;
  wire p14_not_valid;
  wire p13_enable;
  wire p13_data_enable;
  wire p13_not_valid;
  wire p12_enable;
  wire p12_data_enable;
  wire p12_not_valid;
  wire p11_enable;
  wire p11_data_enable;
  wire p11_not_valid;
  wire p10_enable;
  wire p10_data_enable;
  wire p10_not_valid;
  wire p9_enable;
  wire p9_data_enable;
  wire p9_not_valid;
  wire p8_enable;
  wire p8_data_enable;
  wire p8_not_valid;
  wire p7_enable;
  wire p7_data_enable;
  wire p7_not_valid;
  wire p6_enable;
  wire p6_data_enable;
  wire p6_not_valid;
  wire p5_enable;
  wire p5_data_enable;
  wire p5_not_valid;
  wire p4_enable;
  wire p4_data_enable;
  wire p4_not_valid;
  wire p3_enable;
  wire p3_data_enable;
  wire p3_not_valid;
  wire p2_enable;
  wire p2_data_enable;
  wire p2_not_valid;
  wire p1_enable;
  wire [31:0] sub_8463;
  wire [32:0] r__57;
  wire [31:0] concat_8383;
  wire [31:0] r__90;
  wire [31:0] sub_8141;
  wire [32:0] r__47;
  wire [31:0] concat_8061;
  wire [31:0] r__85;
  wire [31:0] sub_7819;
  wire [32:0] r__37;
  wire [31:0] concat_7739;
  wire [31:0] r__80;
  wire [31:0] sub_7497;
  wire [32:0] r__27;
  wire [31:0] concat_7417;
  wire [31:0] r__75;
  wire [31:0] sub_7175;
  wire [32:0] r__17;
  wire [31:0] concat_7095;
  wire [31:0] r__70;
  wire [31:0] sub_6853;
  wire [32:0] r__7;
  wire [31:0] concat_6773;
  wire [31:0] r__65;
  wire p1_data_enable;
  wire p1_not_valid;
  wire [31:0] r__94;
  wire uge_8384;
  wire [31:0] sub_8385;
  wire [32:0] r__55;
  wire [31:0] concat_8303;
  wire [31:0] r__89;
  wire uge_8062;
  wire [31:0] sub_8063;
  wire [32:0] r__45;
  wire [31:0] concat_7981;
  wire [31:0] r__84;
  wire uge_7740;
  wire [31:0] sub_7741;
  wire [32:0] r__35;
  wire [31:0] concat_7659;
  wire [31:0] r__79;
  wire uge_7418;
  wire [31:0] sub_7419;
  wire [32:0] r__25;
  wire [31:0] concat_7337;
  wire [31:0] r__74;
  wire uge_7096;
  wire [31:0] sub_7097;
  wire [32:0] r__15;
  wire [31:0] concat_7015;
  wire [31:0] r__69;
  wire uge_6774;
  wire [31:0] sub_6775;
  wire [32:0] r__5;
  wire [31:0] concat_6693;
  wire p0_enable;
  wire p0_all_active_inputs_valid;
  wire [31:0] r__95;
  wire [31:0] r__93;
  wire uge_8304;
  wire [31:0] sub_8305;
  wire [32:0] r__53;
  wire [31:0] concat_8225;
  wire [31:0] r__88;
  wire uge_7982;
  wire [31:0] sub_7983;
  wire [32:0] r__43;
  wire [31:0] concat_7903;
  wire [31:0] r__83;
  wire uge_7660;
  wire [31:0] sub_7661;
  wire [32:0] r__33;
  wire [31:0] concat_7581;
  wire [31:0] r__78;
  wire uge_7338;
  wire [31:0] sub_7339;
  wire [32:0] r__23;
  wire [31:0] concat_7259;
  wire [31:0] r__73;
  wire uge_7016;
  wire [31:0] sub_7017;
  wire [32:0] r__13;
  wire [31:0] concat_6937;
  wire [31:0] r__68;
  wire uge_6694;
  wire [31:0] sub_6695;
  wire [32:0] r__3;
  wire [32:0] bivisor__1;
  wire [31:0] concat_6615;
  wire p0_data_enable;
  wire lhs_valid_inv;
  wire rhs_valid_inv;
  wire [32:0] r__63;
  wire [32:0] r__61;
  wire [31:0] concat_8467;
  wire [32:0] r__59;
  wire [31:0] r__92;
  wire uge_8226;
  wire [31:0] sub_8227;
  wire [32:0] r__51;
  wire [31:0] concat_8145;
  wire [32:0] r__49;
  wire [31:0] r__87;
  wire uge_7904;
  wire [31:0] sub_7905;
  wire [32:0] r__41;
  wire [31:0] concat_7823;
  wire [32:0] r__39;
  wire [31:0] r__82;
  wire uge_7582;
  wire [31:0] sub_7583;
  wire [32:0] r__31;
  wire [31:0] concat_7501;
  wire [32:0] r__29;
  wire [31:0] r__77;
  wire uge_7260;
  wire [31:0] sub_7261;
  wire [32:0] r__21;
  wire [31:0] concat_7179;
  wire [32:0] r__19;
  wire [31:0] r__72;
  wire uge_6938;
  wire [31:0] sub_6939;
  wire [32:0] r__11;
  wire [31:0] concat_6857;
  wire [32:0] r__9;
  wire [31:0] r__67;
  wire uge_6616;
  wire [31:0] sub_6617;
  wire [31:0] concat_6500;
  wire lhs_valid_load_en;
  wire rhs_valid_load_en;
  wire q__32_squeezed_portion_0_width_1;
  wire p30_enable;
  wire p29_enable;
  wire p28_enable;
  wire p27_enable;
  wire p26_enable;
  wire p25_enable;
  wire uge_8468;
  wire [31:0] sub_8469;
  wire [31:0] concat_8389;
  wire uge_8390;
  wire [30:0] bit_slice_8307;
  wire [31:0] r__91;
  wire uge_8146;
  wire [31:0] sub_8147;
  wire [31:0] concat_8067;
  wire uge_8068;
  wire [30:0] bit_slice_7985;
  wire [31:0] r__86;
  wire uge_7824;
  wire [31:0] sub_7825;
  wire [31:0] concat_7745;
  wire uge_7746;
  wire [30:0] bit_slice_7663;
  wire [31:0] r__81;
  wire uge_7502;
  wire [31:0] sub_7503;
  wire [31:0] concat_7423;
  wire uge_7424;
  wire [30:0] bit_slice_7341;
  wire [31:0] r__76;
  wire uge_7180;
  wire [31:0] sub_7181;
  wire [31:0] concat_7101;
  wire uge_7102;
  wire [30:0] bit_slice_7019;
  wire [31:0] r__71;
  wire uge_6858;
  wire [31:0] sub_6859;
  wire [31:0] concat_6779;
  wire uge_6780;
  wire [30:0] bit_slice_6697;
  wire [31:0] r__66;
  wire uge_6502;
  wire [31:0] sub_6503;
  wire bit_slice_6504;
  wire bit_slice_6505;
  wire bit_slice_6506;
  wire bit_slice_6507;
  wire bit_slice_6508;
  wire bit_slice_6509;
  wire bit_slice_6510;
  wire bit_slice_6511;
  wire bit_slice_6512;
  wire bit_slice_6513;
  wire bit_slice_6514;
  wire bit_slice_6515;
  wire bit_slice_6516;
  wire bit_slice_6517;
  wire bit_slice_6518;
  wire bit_slice_6519;
  wire bit_slice_6520;
  wire bit_slice_6521;
  wire bit_slice_6522;
  wire bit_slice_6523;
  wire bit_slice_6524;
  wire bit_slice_6525;
  wire bit_slice_6526;
  wire bit_slice_6527;
  wire bit_slice_6528;
  wire bit_slice_6529;
  wire bit_slice_6530;
  wire bit_slice_6531;
  wire bit_slice_6532;
  wire bit_slice_6533;
  wire bit_slice_6534;
  wire lhs_load_en;
  wire rhs_load_en;
  wire [31:0] q__32;
  assign result_valid_inv = ~result_valid_reg;
  assign result_valid_load_en = result_ready | result_valid_inv;
  assign result_load_en = p24_valid & result_valid_load_en;
  assign p25_stage_done = p24_valid & result_load_en;
  assign p25_not_valid = ~p24_valid;
  assign p24_enable = p25_stage_done | p25_not_valid;
  assign p24_data_enable = p24_enable & p23_valid;
  assign p24_not_valid = ~p23_valid;
  assign p23_enable = p24_data_enable | p24_not_valid;
  assign p23_data_enable = p23_enable & p22_valid;
  assign p23_not_valid = ~p22_valid;
  assign p22_enable = p23_data_enable | p23_not_valid;
  assign p22_data_enable = p22_enable & p21_valid;
  assign p22_not_valid = ~p21_valid;
  assign p21_enable = p22_data_enable | p22_not_valid;
  assign p21_data_enable = p21_enable & p20_valid;
  assign p21_not_valid = ~p20_valid;
  assign p20_enable = p21_data_enable | p21_not_valid;
  assign p20_data_enable = p20_enable & p19_valid;
  assign p20_not_valid = ~p19_valid;
  assign p19_enable = p20_data_enable | p20_not_valid;
  assign p19_data_enable = p19_enable & p18_valid;
  assign p19_not_valid = ~p18_valid;
  assign p18_enable = p19_data_enable | p19_not_valid;
  assign p18_data_enable = p18_enable & p17_valid;
  assign p18_not_valid = ~p17_valid;
  assign p17_enable = p18_data_enable | p18_not_valid;
  assign p17_data_enable = p17_enable & p16_valid;
  assign p17_not_valid = ~p16_valid;
  assign p16_enable = p17_data_enable | p17_not_valid;
  assign p16_data_enable = p16_enable & p15_valid;
  assign p16_not_valid = ~p15_valid;
  assign p15_enable = p16_data_enable | p16_not_valid;
  assign p15_data_enable = p15_enable & p14_valid;
  assign p15_not_valid = ~p14_valid;
  assign p14_enable = p15_data_enable | p15_not_valid;
  assign p14_data_enable = p14_enable & p13_valid;
  assign p14_not_valid = ~p13_valid;
  assign p13_enable = p14_data_enable | p14_not_valid;
  assign p13_data_enable = p13_enable & p12_valid;
  assign p13_not_valid = ~p12_valid;
  assign p12_enable = p13_data_enable | p13_not_valid;
  assign p12_data_enable = p12_enable & p11_valid;
  assign p12_not_valid = ~p11_valid;
  assign p11_enable = p12_data_enable | p12_not_valid;
  assign p11_data_enable = p11_enable & p10_valid;
  assign p11_not_valid = ~p10_valid;
  assign p10_enable = p11_data_enable | p11_not_valid;
  assign p10_data_enable = p10_enable & p9_valid;
  assign p10_not_valid = ~p9_valid;
  assign p9_enable = p10_data_enable | p10_not_valid;
  assign p9_data_enable = p9_enable & p8_valid;
  assign p9_not_valid = ~p8_valid;
  assign p8_enable = p9_data_enable | p9_not_valid;
  assign p8_data_enable = p8_enable & p7_valid;
  assign p8_not_valid = ~p7_valid;
  assign p7_enable = p8_data_enable | p8_not_valid;
  assign p7_data_enable = p7_enable & p6_valid;
  assign p7_not_valid = ~p6_valid;
  assign p6_enable = p7_data_enable | p7_not_valid;
  assign p6_data_enable = p6_enable & p5_valid;
  assign p6_not_valid = ~p5_valid;
  assign p5_enable = p6_data_enable | p6_not_valid;
  assign p5_data_enable = p5_enable & p4_valid;
  assign p5_not_valid = ~p4_valid;
  assign p4_enable = p5_data_enable | p5_not_valid;
  assign p4_data_enable = p4_enable & p3_valid;
  assign p4_not_valid = ~p3_valid;
  assign p3_enable = p4_data_enable | p4_not_valid;
  assign p3_data_enable = p3_enable & p2_valid;
  assign p3_not_valid = ~p2_valid;
  assign p2_enable = p3_data_enable | p3_not_valid;
  assign p2_data_enable = p2_enable & p1_valid;
  assign p2_not_valid = ~p1_valid;
  assign p1_enable = p2_data_enable | p2_not_valid;
  assign sub_8463 = p23_concat_8389 - p23_b;
  assign r__57 = {p22_r__92, p22_bit_slice_6531};
  assign concat_8383 = {p22_bit_slice_8307, p22_bit_slice_6531};
  assign r__90 = p20_uge_8146 ? p20_sub_8147 : p20_concat_8145;
  assign sub_8141 = p19_concat_8067 - p19_b;
  assign r__47 = {p18_r__87, p18_bit_slice_6526};
  assign concat_8061 = {p18_bit_slice_7985, p18_bit_slice_6526};
  assign r__85 = p16_uge_7824 ? p16_sub_7825 : p16_concat_7823;
  assign sub_7819 = p15_concat_7745 - p15_b;
  assign r__37 = {p14_r__82, p14_bit_slice_6521};
  assign concat_7739 = {p14_bit_slice_7663, p14_bit_slice_6521};
  assign r__80 = p12_uge_7502 ? p12_sub_7503 : p12_concat_7501;
  assign sub_7497 = p11_concat_7423 - p11_b;
  assign r__27 = {p10_r__77, p10_bit_slice_6516};
  assign concat_7417 = {p10_bit_slice_7341, p10_bit_slice_6516};
  assign r__75 = p8_uge_7180 ? p8_sub_7181 : p8_concat_7179;
  assign sub_7175 = p7_concat_7101 - p7_b;
  assign r__17 = {p6_r__72, p6_bit_slice_6511};
  assign concat_7095 = {p6_bit_slice_7019, p6_bit_slice_6511};
  assign r__70 = p4_uge_6858 ? p4_sub_6859 : p4_concat_6857;
  assign sub_6853 = p3_concat_6779 - p3_b;
  assign r__7 = {p2_r__67, p2_bit_slice_6506};
  assign concat_6773 = {p2_bit_slice_6697, p2_bit_slice_6506};
  assign r__65 = p0_uge_6502 ? p0_sub_6503 : p0_concat_6500;
  assign p1_data_enable = p1_enable & p0_valid;
  assign p1_not_valid = ~p0_valid;
  assign r__94 = p23_uge_8390 ? sub_8463 : p23_concat_8389;
  assign uge_8384 = r__57 >= p22_bivisor__1;
  assign sub_8385 = concat_8383 - p22_b;
  assign r__55 = {p21_r__91, p21_bit_slice_6530};
  assign concat_8303 = {p21_r__91[30:0], p21_bit_slice_6530};
  assign r__89 = p19_uge_8068 ? sub_8141 : p19_concat_8067;
  assign uge_8062 = r__47 >= p18_bivisor__1;
  assign sub_8063 = concat_8061 - p18_b;
  assign r__45 = {p17_r__86, p17_bit_slice_6525};
  assign concat_7981 = {p17_r__86[30:0], p17_bit_slice_6525};
  assign r__84 = p15_uge_7746 ? sub_7819 : p15_concat_7745;
  assign uge_7740 = r__37 >= p14_bivisor__1;
  assign sub_7741 = concat_7739 - p14_b;
  assign r__35 = {p13_r__81, p13_bit_slice_6520};
  assign concat_7659 = {p13_r__81[30:0], p13_bit_slice_6520};
  assign r__79 = p11_uge_7424 ? sub_7497 : p11_concat_7423;
  assign uge_7418 = r__27 >= p10_bivisor__1;
  assign sub_7419 = concat_7417 - p10_b;
  assign r__25 = {p9_r__76, p9_bit_slice_6515};
  assign concat_7337 = {p9_r__76[30:0], p9_bit_slice_6515};
  assign r__74 = p7_uge_7102 ? sub_7175 : p7_concat_7101;
  assign uge_7096 = r__17 >= p6_bivisor__1;
  assign sub_7097 = concat_7095 - p6_b;
  assign r__15 = {p5_r__71, p5_bit_slice_6510};
  assign concat_7015 = {p5_r__71[30:0], p5_bit_slice_6510};
  assign r__69 = p3_uge_6780 ? sub_6853 : p3_concat_6779;
  assign uge_6774 = r__7 >= p2_bivisor__1;
  assign sub_6775 = concat_6773 - p2_b;
  assign r__5 = {p1_r__66, p1_bit_slice_6505};
  assign concat_6693 = {p1_r__66[30:0], p1_bit_slice_6505};
  assign p0_enable = p1_data_enable | p1_not_valid;
  assign p0_all_active_inputs_valid = lhs_valid_reg & rhs_valid_reg;
  assign r__95 = p24_uge_8468 ? p24_sub_8469 : p24_concat_8467;
  assign r__93 = uge_8384 ? sub_8385 : concat_8383;
  assign uge_8304 = r__55 >= p21_bivisor__1;
  assign sub_8305 = concat_8303 - p21_b;
  assign r__53 = {r__90, p20_bit_slice_6529};
  assign concat_8225 = {r__90[30:0], p20_bit_slice_6529};
  assign r__88 = uge_8062 ? sub_8063 : concat_8061;
  assign uge_7982 = r__45 >= p17_bivisor__1;
  assign sub_7983 = concat_7981 - p17_b;
  assign r__43 = {r__85, p16_bit_slice_6524};
  assign concat_7903 = {r__85[30:0], p16_bit_slice_6524};
  assign r__83 = uge_7740 ? sub_7741 : concat_7739;
  assign uge_7660 = r__35 >= p13_bivisor__1;
  assign sub_7661 = concat_7659 - p13_b;
  assign r__33 = {r__80, p12_bit_slice_6519};
  assign concat_7581 = {r__80[30:0], p12_bit_slice_6519};
  assign r__78 = uge_7418 ? sub_7419 : concat_7417;
  assign uge_7338 = r__25 >= p9_bivisor__1;
  assign sub_7339 = concat_7337 - p9_b;
  assign r__23 = {r__75, p8_bit_slice_6514};
  assign concat_7259 = {r__75[30:0], p8_bit_slice_6514};
  assign r__73 = uge_7096 ? sub_7097 : concat_7095;
  assign uge_7016 = r__15 >= p5_bivisor__1;
  assign sub_7017 = concat_7015 - p5_b;
  assign r__13 = {r__70, p4_bit_slice_6509};
  assign concat_6937 = {r__70[30:0], p4_bit_slice_6509};
  assign r__68 = uge_6774 ? sub_6775 : concat_6773;
  assign uge_6694 = r__5 >= p1_bivisor__1;
  assign sub_6695 = concat_6693 - p1_b;
  assign r__3 = {r__65, p0_bit_slice_6504};
  assign bivisor__1 = {1'h0, p0_b};
  assign concat_6615 = {r__65[30:0], p0_bit_slice_6504};
  assign p0_data_enable = p0_enable & p0_all_active_inputs_valid;
  assign lhs_valid_inv = ~lhs_valid_reg;
  assign rhs_valid_inv = ~rhs_valid_reg;
  assign r__63 = {r__95, p24_bit_slice_6534};
  assign r__61 = {r__94, p23_bit_slice_6533};
  assign concat_8467 = {r__94[30:0], p23_bit_slice_6533};
  assign r__59 = {r__93, p22_bit_slice_6532};
  assign r__92 = uge_8304 ? sub_8305 : concat_8303;
  assign uge_8226 = r__53 >= p20_bivisor__1;
  assign sub_8227 = concat_8225 - p20_b;
  assign r__51 = {r__89, p19_bit_slice_6528};
  assign concat_8145 = {r__89[30:0], p19_bit_slice_6528};
  assign r__49 = {r__88, p18_bit_slice_6527};
  assign r__87 = uge_7982 ? sub_7983 : concat_7981;
  assign uge_7904 = r__43 >= p16_bivisor__1;
  assign sub_7905 = concat_7903 - p16_b;
  assign r__41 = {r__84, p15_bit_slice_6523};
  assign concat_7823 = {r__84[30:0], p15_bit_slice_6523};
  assign r__39 = {r__83, p14_bit_slice_6522};
  assign r__82 = uge_7660 ? sub_7661 : concat_7659;
  assign uge_7582 = r__33 >= p12_bivisor__1;
  assign sub_7583 = concat_7581 - p12_b;
  assign r__31 = {r__79, p11_bit_slice_6518};
  assign concat_7501 = {r__79[30:0], p11_bit_slice_6518};
  assign r__29 = {r__78, p10_bit_slice_6517};
  assign r__77 = uge_7338 ? sub_7339 : concat_7337;
  assign uge_7260 = r__23 >= p8_bivisor__1;
  assign sub_7261 = concat_7259 - p8_b;
  assign r__21 = {r__74, p7_bit_slice_6513};
  assign concat_7179 = {r__74[30:0], p7_bit_slice_6513};
  assign r__19 = {r__73, p6_bit_slice_6512};
  assign r__72 = uge_7016 ? sub_7017 : concat_7015;
  assign uge_6938 = r__13 >= p4_bivisor__1;
  assign sub_6939 = concat_6937 - p4_b;
  assign r__11 = {r__69, p3_bit_slice_6508};
  assign concat_6857 = {r__69[30:0], p3_bit_slice_6508};
  assign r__9 = {r__68, p2_bit_slice_6507};
  assign r__67 = uge_6694 ? sub_6695 : concat_6693;
  assign uge_6616 = r__3 >= bivisor__1;
  assign sub_6617 = concat_6615 - p0_b;
  assign concat_6500 = {31'h0000_0000, lhs_reg[31]};
  assign lhs_valid_load_en = p0_data_enable | lhs_valid_inv;
  assign rhs_valid_load_en = p0_data_enable | rhs_valid_inv;
  assign q__32_squeezed_portion_0_width_1 = r__63 >= p24_bivisor__1;
  assign p30_enable = 1'h1;
  assign p29_enable = 1'h1;
  assign p28_enable = 1'h1;
  assign p27_enable = 1'h1;
  assign p26_enable = 1'h1;
  assign p25_enable = 1'h1;
  assign uge_8468 = r__61 >= p23_bivisor__1;
  assign sub_8469 = concat_8467 - p23_b;
  assign concat_8389 = {r__93[30:0], p22_bit_slice_6532};
  assign uge_8390 = r__59 >= p22_bivisor__1;
  assign bit_slice_8307 = r__92[30:0];
  assign r__91 = uge_8226 ? sub_8227 : concat_8225;
  assign uge_8146 = r__51 >= p19_bivisor__1;
  assign sub_8147 = concat_8145 - p19_b;
  assign concat_8067 = {r__88[30:0], p18_bit_slice_6527};
  assign uge_8068 = r__49 >= p18_bivisor__1;
  assign bit_slice_7985 = r__87[30:0];
  assign r__86 = uge_7904 ? sub_7905 : concat_7903;
  assign uge_7824 = r__41 >= p15_bivisor__1;
  assign sub_7825 = concat_7823 - p15_b;
  assign concat_7745 = {r__83[30:0], p14_bit_slice_6522};
  assign uge_7746 = r__39 >= p14_bivisor__1;
  assign bit_slice_7663 = r__82[30:0];
  assign r__81 = uge_7582 ? sub_7583 : concat_7581;
  assign uge_7502 = r__31 >= p11_bivisor__1;
  assign sub_7503 = concat_7501 - p11_b;
  assign concat_7423 = {r__78[30:0], p10_bit_slice_6517};
  assign uge_7424 = r__29 >= p10_bivisor__1;
  assign bit_slice_7341 = r__77[30:0];
  assign r__76 = uge_7260 ? sub_7261 : concat_7259;
  assign uge_7180 = r__21 >= p7_bivisor__1;
  assign sub_7181 = concat_7179 - p7_b;
  assign concat_7101 = {r__73[30:0], p6_bit_slice_6512};
  assign uge_7102 = r__19 >= p6_bivisor__1;
  assign bit_slice_7019 = r__72[30:0];
  assign r__71 = uge_6938 ? sub_6939 : concat_6937;
  assign uge_6858 = r__11 >= p3_bivisor__1;
  assign sub_6859 = concat_6857 - p3_b;
  assign concat_6779 = {r__68[30:0], p2_bit_slice_6507};
  assign uge_6780 = r__9 >= p2_bivisor__1;
  assign bit_slice_6697 = r__67[30:0];
  assign r__66 = uge_6616 ? sub_6617 : concat_6615;
  assign uge_6502 = concat_6500 >= rhs_reg;
  assign sub_6503 = concat_6500 - rhs_reg;
  assign bit_slice_6504 = lhs_reg[30];
  assign bit_slice_6505 = lhs_reg[29];
  assign bit_slice_6506 = lhs_reg[28];
  assign bit_slice_6507 = lhs_reg[27];
  assign bit_slice_6508 = lhs_reg[26];
  assign bit_slice_6509 = lhs_reg[25];
  assign bit_slice_6510 = lhs_reg[24];
  assign bit_slice_6511 = lhs_reg[23];
  assign bit_slice_6512 = lhs_reg[22];
  assign bit_slice_6513 = lhs_reg[21];
  assign bit_slice_6514 = lhs_reg[20];
  assign bit_slice_6515 = lhs_reg[19];
  assign bit_slice_6516 = lhs_reg[18];
  assign bit_slice_6517 = lhs_reg[17];
  assign bit_slice_6518 = lhs_reg[16];
  assign bit_slice_6519 = lhs_reg[15];
  assign bit_slice_6520 = lhs_reg[14];
  assign bit_slice_6521 = lhs_reg[13];
  assign bit_slice_6522 = lhs_reg[12];
  assign bit_slice_6523 = lhs_reg[11];
  assign bit_slice_6524 = lhs_reg[10];
  assign bit_slice_6525 = lhs_reg[9];
  assign bit_slice_6526 = lhs_reg[8];
  assign bit_slice_6527 = lhs_reg[7];
  assign bit_slice_6528 = lhs_reg[6];
  assign bit_slice_6529 = lhs_reg[5];
  assign bit_slice_6530 = lhs_reg[4];
  assign bit_slice_6531 = lhs_reg[3];
  assign bit_slice_6532 = lhs_reg[2];
  assign bit_slice_6533 = lhs_reg[1];
  assign bit_slice_6534 = lhs_reg[0];
  assign lhs_load_en = lhs_valid & lhs_valid_load_en;
  assign rhs_load_en = rhs_valid & rhs_valid_load_en;
  assign q__32 = {p24_uge_6502, p24_uge_6616, p24_uge_6694, p24_uge_6774, p24_uge_6780, p24_uge_6858, p24_uge_6938, p24_uge_7016, p24_uge_7096, p24_uge_7102, p24_uge_7180, p24_uge_7260, p24_uge_7338, p24_uge_7418, p24_uge_7424, p24_uge_7502, p24_uge_7582, p24_uge_7660, p24_uge_7740, p24_uge_7746, p24_uge_7824, p24_uge_7904, p24_uge_7982, p24_uge_8062, p24_uge_8068, p24_uge_8146, p24_uge_8226, p24_uge_8304, p24_uge_8384, p24_uge_8390, p24_uge_8468, q__32_squeezed_portion_0_width_1};
  always @ (posedge clk) begin
    if (rst) begin
      p0_concat_6500 <= 32'h0000_0000;
      p0_b <= 32'h0000_0000;
      p0_uge_6502 <= 1'h0;
      p0_sub_6503 <= 32'h0000_0000;
      p0_bit_slice_6504 <= 1'h0;
      p0_bit_slice_6505 <= 1'h0;
      p0_bit_slice_6506 <= 1'h0;
      p0_bit_slice_6507 <= 1'h0;
      p0_bit_slice_6508 <= 1'h0;
      p0_bit_slice_6509 <= 1'h0;
      p0_bit_slice_6510 <= 1'h0;
      p0_bit_slice_6511 <= 1'h0;
      p0_bit_slice_6512 <= 1'h0;
      p0_bit_slice_6513 <= 1'h0;
      p0_bit_slice_6514 <= 1'h0;
      p0_bit_slice_6515 <= 1'h0;
      p0_bit_slice_6516 <= 1'h0;
      p0_bit_slice_6517 <= 1'h0;
      p0_bit_slice_6518 <= 1'h0;
      p0_bit_slice_6519 <= 1'h0;
      p0_bit_slice_6520 <= 1'h0;
      p0_bit_slice_6521 <= 1'h0;
      p0_bit_slice_6522 <= 1'h0;
      p0_bit_slice_6523 <= 1'h0;
      p0_bit_slice_6524 <= 1'h0;
      p0_bit_slice_6525 <= 1'h0;
      p0_bit_slice_6526 <= 1'h0;
      p0_bit_slice_6527 <= 1'h0;
      p0_bit_slice_6528 <= 1'h0;
      p0_bit_slice_6529 <= 1'h0;
      p0_bit_slice_6530 <= 1'h0;
      p0_bit_slice_6531 <= 1'h0;
      p0_bit_slice_6532 <= 1'h0;
      p0_bit_slice_6533 <= 1'h0;
      p0_bit_slice_6534 <= 1'h0;
      p1_b <= 32'h0000_0000;
      p1_uge_6502 <= 1'h0;
      p1_bivisor__1 <= 33'h0_0000_0000;
      p1_uge_6616 <= 1'h0;
      p1_r__66 <= 32'h0000_0000;
      p1_bit_slice_6505 <= 1'h0;
      p1_bit_slice_6506 <= 1'h0;
      p1_bit_slice_6507 <= 1'h0;
      p1_bit_slice_6508 <= 1'h0;
      p1_bit_slice_6509 <= 1'h0;
      p1_bit_slice_6510 <= 1'h0;
      p1_bit_slice_6511 <= 1'h0;
      p1_bit_slice_6512 <= 1'h0;
      p1_bit_slice_6513 <= 1'h0;
      p1_bit_slice_6514 <= 1'h0;
      p1_bit_slice_6515 <= 1'h0;
      p1_bit_slice_6516 <= 1'h0;
      p1_bit_slice_6517 <= 1'h0;
      p1_bit_slice_6518 <= 1'h0;
      p1_bit_slice_6519 <= 1'h0;
      p1_bit_slice_6520 <= 1'h0;
      p1_bit_slice_6521 <= 1'h0;
      p1_bit_slice_6522 <= 1'h0;
      p1_bit_slice_6523 <= 1'h0;
      p1_bit_slice_6524 <= 1'h0;
      p1_bit_slice_6525 <= 1'h0;
      p1_bit_slice_6526 <= 1'h0;
      p1_bit_slice_6527 <= 1'h0;
      p1_bit_slice_6528 <= 1'h0;
      p1_bit_slice_6529 <= 1'h0;
      p1_bit_slice_6530 <= 1'h0;
      p1_bit_slice_6531 <= 1'h0;
      p1_bit_slice_6532 <= 1'h0;
      p1_bit_slice_6533 <= 1'h0;
      p1_bit_slice_6534 <= 1'h0;
      p2_b <= 32'h0000_0000;
      p2_uge_6502 <= 1'h0;
      p2_bivisor__1 <= 33'h0_0000_0000;
      p2_uge_6616 <= 1'h0;
      p2_uge_6694 <= 1'h0;
      p2_r__67 <= 32'h0000_0000;
      p2_bit_slice_6506 <= 1'h0;
      p2_bit_slice_6697 <= 31'h0000_0000;
      p2_bit_slice_6507 <= 1'h0;
      p2_bit_slice_6508 <= 1'h0;
      p2_bit_slice_6509 <= 1'h0;
      p2_bit_slice_6510 <= 1'h0;
      p2_bit_slice_6511 <= 1'h0;
      p2_bit_slice_6512 <= 1'h0;
      p2_bit_slice_6513 <= 1'h0;
      p2_bit_slice_6514 <= 1'h0;
      p2_bit_slice_6515 <= 1'h0;
      p2_bit_slice_6516 <= 1'h0;
      p2_bit_slice_6517 <= 1'h0;
      p2_bit_slice_6518 <= 1'h0;
      p2_bit_slice_6519 <= 1'h0;
      p2_bit_slice_6520 <= 1'h0;
      p2_bit_slice_6521 <= 1'h0;
      p2_bit_slice_6522 <= 1'h0;
      p2_bit_slice_6523 <= 1'h0;
      p2_bit_slice_6524 <= 1'h0;
      p2_bit_slice_6525 <= 1'h0;
      p2_bit_slice_6526 <= 1'h0;
      p2_bit_slice_6527 <= 1'h0;
      p2_bit_slice_6528 <= 1'h0;
      p2_bit_slice_6529 <= 1'h0;
      p2_bit_slice_6530 <= 1'h0;
      p2_bit_slice_6531 <= 1'h0;
      p2_bit_slice_6532 <= 1'h0;
      p2_bit_slice_6533 <= 1'h0;
      p2_bit_slice_6534 <= 1'h0;
      p3_b <= 32'h0000_0000;
      p3_uge_6502 <= 1'h0;
      p3_bivisor__1 <= 33'h0_0000_0000;
      p3_uge_6616 <= 1'h0;
      p3_uge_6694 <= 1'h0;
      p3_uge_6774 <= 1'h0;
      p3_concat_6779 <= 32'h0000_0000;
      p3_uge_6780 <= 1'h0;
      p3_bit_slice_6508 <= 1'h0;
      p3_bit_slice_6509 <= 1'h0;
      p3_bit_slice_6510 <= 1'h0;
      p3_bit_slice_6511 <= 1'h0;
      p3_bit_slice_6512 <= 1'h0;
      p3_bit_slice_6513 <= 1'h0;
      p3_bit_slice_6514 <= 1'h0;
      p3_bit_slice_6515 <= 1'h0;
      p3_bit_slice_6516 <= 1'h0;
      p3_bit_slice_6517 <= 1'h0;
      p3_bit_slice_6518 <= 1'h0;
      p3_bit_slice_6519 <= 1'h0;
      p3_bit_slice_6520 <= 1'h0;
      p3_bit_slice_6521 <= 1'h0;
      p3_bit_slice_6522 <= 1'h0;
      p3_bit_slice_6523 <= 1'h0;
      p3_bit_slice_6524 <= 1'h0;
      p3_bit_slice_6525 <= 1'h0;
      p3_bit_slice_6526 <= 1'h0;
      p3_bit_slice_6527 <= 1'h0;
      p3_bit_slice_6528 <= 1'h0;
      p3_bit_slice_6529 <= 1'h0;
      p3_bit_slice_6530 <= 1'h0;
      p3_bit_slice_6531 <= 1'h0;
      p3_bit_slice_6532 <= 1'h0;
      p3_bit_slice_6533 <= 1'h0;
      p3_bit_slice_6534 <= 1'h0;
      p4_b <= 32'h0000_0000;
      p4_uge_6502 <= 1'h0;
      p4_bivisor__1 <= 33'h0_0000_0000;
      p4_uge_6616 <= 1'h0;
      p4_uge_6694 <= 1'h0;
      p4_uge_6774 <= 1'h0;
      p4_uge_6780 <= 1'h0;
      p4_concat_6857 <= 32'h0000_0000;
      p4_uge_6858 <= 1'h0;
      p4_sub_6859 <= 32'h0000_0000;
      p4_bit_slice_6509 <= 1'h0;
      p4_bit_slice_6510 <= 1'h0;
      p4_bit_slice_6511 <= 1'h0;
      p4_bit_slice_6512 <= 1'h0;
      p4_bit_slice_6513 <= 1'h0;
      p4_bit_slice_6514 <= 1'h0;
      p4_bit_slice_6515 <= 1'h0;
      p4_bit_slice_6516 <= 1'h0;
      p4_bit_slice_6517 <= 1'h0;
      p4_bit_slice_6518 <= 1'h0;
      p4_bit_slice_6519 <= 1'h0;
      p4_bit_slice_6520 <= 1'h0;
      p4_bit_slice_6521 <= 1'h0;
      p4_bit_slice_6522 <= 1'h0;
      p4_bit_slice_6523 <= 1'h0;
      p4_bit_slice_6524 <= 1'h0;
      p4_bit_slice_6525 <= 1'h0;
      p4_bit_slice_6526 <= 1'h0;
      p4_bit_slice_6527 <= 1'h0;
      p4_bit_slice_6528 <= 1'h0;
      p4_bit_slice_6529 <= 1'h0;
      p4_bit_slice_6530 <= 1'h0;
      p4_bit_slice_6531 <= 1'h0;
      p4_bit_slice_6532 <= 1'h0;
      p4_bit_slice_6533 <= 1'h0;
      p4_bit_slice_6534 <= 1'h0;
      p5_b <= 32'h0000_0000;
      p5_uge_6502 <= 1'h0;
      p5_bivisor__1 <= 33'h0_0000_0000;
      p5_uge_6616 <= 1'h0;
      p5_uge_6694 <= 1'h0;
      p5_uge_6774 <= 1'h0;
      p5_uge_6780 <= 1'h0;
      p5_uge_6858 <= 1'h0;
      p5_uge_6938 <= 1'h0;
      p5_r__71 <= 32'h0000_0000;
      p5_bit_slice_6510 <= 1'h0;
      p5_bit_slice_6511 <= 1'h0;
      p5_bit_slice_6512 <= 1'h0;
      p5_bit_slice_6513 <= 1'h0;
      p5_bit_slice_6514 <= 1'h0;
      p5_bit_slice_6515 <= 1'h0;
      p5_bit_slice_6516 <= 1'h0;
      p5_bit_slice_6517 <= 1'h0;
      p5_bit_slice_6518 <= 1'h0;
      p5_bit_slice_6519 <= 1'h0;
      p5_bit_slice_6520 <= 1'h0;
      p5_bit_slice_6521 <= 1'h0;
      p5_bit_slice_6522 <= 1'h0;
      p5_bit_slice_6523 <= 1'h0;
      p5_bit_slice_6524 <= 1'h0;
      p5_bit_slice_6525 <= 1'h0;
      p5_bit_slice_6526 <= 1'h0;
      p5_bit_slice_6527 <= 1'h0;
      p5_bit_slice_6528 <= 1'h0;
      p5_bit_slice_6529 <= 1'h0;
      p5_bit_slice_6530 <= 1'h0;
      p5_bit_slice_6531 <= 1'h0;
      p5_bit_slice_6532 <= 1'h0;
      p5_bit_slice_6533 <= 1'h0;
      p5_bit_slice_6534 <= 1'h0;
      p6_b <= 32'h0000_0000;
      p6_uge_6502 <= 1'h0;
      p6_bivisor__1 <= 33'h0_0000_0000;
      p6_uge_6616 <= 1'h0;
      p6_uge_6694 <= 1'h0;
      p6_uge_6774 <= 1'h0;
      p6_uge_6780 <= 1'h0;
      p6_uge_6858 <= 1'h0;
      p6_uge_6938 <= 1'h0;
      p6_uge_7016 <= 1'h0;
      p6_r__72 <= 32'h0000_0000;
      p6_bit_slice_6511 <= 1'h0;
      p6_bit_slice_7019 <= 31'h0000_0000;
      p6_bit_slice_6512 <= 1'h0;
      p6_bit_slice_6513 <= 1'h0;
      p6_bit_slice_6514 <= 1'h0;
      p6_bit_slice_6515 <= 1'h0;
      p6_bit_slice_6516 <= 1'h0;
      p6_bit_slice_6517 <= 1'h0;
      p6_bit_slice_6518 <= 1'h0;
      p6_bit_slice_6519 <= 1'h0;
      p6_bit_slice_6520 <= 1'h0;
      p6_bit_slice_6521 <= 1'h0;
      p6_bit_slice_6522 <= 1'h0;
      p6_bit_slice_6523 <= 1'h0;
      p6_bit_slice_6524 <= 1'h0;
      p6_bit_slice_6525 <= 1'h0;
      p6_bit_slice_6526 <= 1'h0;
      p6_bit_slice_6527 <= 1'h0;
      p6_bit_slice_6528 <= 1'h0;
      p6_bit_slice_6529 <= 1'h0;
      p6_bit_slice_6530 <= 1'h0;
      p6_bit_slice_6531 <= 1'h0;
      p6_bit_slice_6532 <= 1'h0;
      p6_bit_slice_6533 <= 1'h0;
      p6_bit_slice_6534 <= 1'h0;
      p7_b <= 32'h0000_0000;
      p7_uge_6502 <= 1'h0;
      p7_bivisor__1 <= 33'h0_0000_0000;
      p7_uge_6616 <= 1'h0;
      p7_uge_6694 <= 1'h0;
      p7_uge_6774 <= 1'h0;
      p7_uge_6780 <= 1'h0;
      p7_uge_6858 <= 1'h0;
      p7_uge_6938 <= 1'h0;
      p7_uge_7016 <= 1'h0;
      p7_uge_7096 <= 1'h0;
      p7_concat_7101 <= 32'h0000_0000;
      p7_uge_7102 <= 1'h0;
      p7_bit_slice_6513 <= 1'h0;
      p7_bit_slice_6514 <= 1'h0;
      p7_bit_slice_6515 <= 1'h0;
      p7_bit_slice_6516 <= 1'h0;
      p7_bit_slice_6517 <= 1'h0;
      p7_bit_slice_6518 <= 1'h0;
      p7_bit_slice_6519 <= 1'h0;
      p7_bit_slice_6520 <= 1'h0;
      p7_bit_slice_6521 <= 1'h0;
      p7_bit_slice_6522 <= 1'h0;
      p7_bit_slice_6523 <= 1'h0;
      p7_bit_slice_6524 <= 1'h0;
      p7_bit_slice_6525 <= 1'h0;
      p7_bit_slice_6526 <= 1'h0;
      p7_bit_slice_6527 <= 1'h0;
      p7_bit_slice_6528 <= 1'h0;
      p7_bit_slice_6529 <= 1'h0;
      p7_bit_slice_6530 <= 1'h0;
      p7_bit_slice_6531 <= 1'h0;
      p7_bit_slice_6532 <= 1'h0;
      p7_bit_slice_6533 <= 1'h0;
      p7_bit_slice_6534 <= 1'h0;
      p8_b <= 32'h0000_0000;
      p8_uge_6502 <= 1'h0;
      p8_bivisor__1 <= 33'h0_0000_0000;
      p8_uge_6616 <= 1'h0;
      p8_uge_6694 <= 1'h0;
      p8_uge_6774 <= 1'h0;
      p8_uge_6780 <= 1'h0;
      p8_uge_6858 <= 1'h0;
      p8_uge_6938 <= 1'h0;
      p8_uge_7016 <= 1'h0;
      p8_uge_7096 <= 1'h0;
      p8_uge_7102 <= 1'h0;
      p8_concat_7179 <= 32'h0000_0000;
      p8_uge_7180 <= 1'h0;
      p8_sub_7181 <= 32'h0000_0000;
      p8_bit_slice_6514 <= 1'h0;
      p8_bit_slice_6515 <= 1'h0;
      p8_bit_slice_6516 <= 1'h0;
      p8_bit_slice_6517 <= 1'h0;
      p8_bit_slice_6518 <= 1'h0;
      p8_bit_slice_6519 <= 1'h0;
      p8_bit_slice_6520 <= 1'h0;
      p8_bit_slice_6521 <= 1'h0;
      p8_bit_slice_6522 <= 1'h0;
      p8_bit_slice_6523 <= 1'h0;
      p8_bit_slice_6524 <= 1'h0;
      p8_bit_slice_6525 <= 1'h0;
      p8_bit_slice_6526 <= 1'h0;
      p8_bit_slice_6527 <= 1'h0;
      p8_bit_slice_6528 <= 1'h0;
      p8_bit_slice_6529 <= 1'h0;
      p8_bit_slice_6530 <= 1'h0;
      p8_bit_slice_6531 <= 1'h0;
      p8_bit_slice_6532 <= 1'h0;
      p8_bit_slice_6533 <= 1'h0;
      p8_bit_slice_6534 <= 1'h0;
      p9_b <= 32'h0000_0000;
      p9_uge_6502 <= 1'h0;
      p9_bivisor__1 <= 33'h0_0000_0000;
      p9_uge_6616 <= 1'h0;
      p9_uge_6694 <= 1'h0;
      p9_uge_6774 <= 1'h0;
      p9_uge_6780 <= 1'h0;
      p9_uge_6858 <= 1'h0;
      p9_uge_6938 <= 1'h0;
      p9_uge_7016 <= 1'h0;
      p9_uge_7096 <= 1'h0;
      p9_uge_7102 <= 1'h0;
      p9_uge_7180 <= 1'h0;
      p9_uge_7260 <= 1'h0;
      p9_r__76 <= 32'h0000_0000;
      p9_bit_slice_6515 <= 1'h0;
      p9_bit_slice_6516 <= 1'h0;
      p9_bit_slice_6517 <= 1'h0;
      p9_bit_slice_6518 <= 1'h0;
      p9_bit_slice_6519 <= 1'h0;
      p9_bit_slice_6520 <= 1'h0;
      p9_bit_slice_6521 <= 1'h0;
      p9_bit_slice_6522 <= 1'h0;
      p9_bit_slice_6523 <= 1'h0;
      p9_bit_slice_6524 <= 1'h0;
      p9_bit_slice_6525 <= 1'h0;
      p9_bit_slice_6526 <= 1'h0;
      p9_bit_slice_6527 <= 1'h0;
      p9_bit_slice_6528 <= 1'h0;
      p9_bit_slice_6529 <= 1'h0;
      p9_bit_slice_6530 <= 1'h0;
      p9_bit_slice_6531 <= 1'h0;
      p9_bit_slice_6532 <= 1'h0;
      p9_bit_slice_6533 <= 1'h0;
      p9_bit_slice_6534 <= 1'h0;
      p10_b <= 32'h0000_0000;
      p10_uge_6502 <= 1'h0;
      p10_bivisor__1 <= 33'h0_0000_0000;
      p10_uge_6616 <= 1'h0;
      p10_uge_6694 <= 1'h0;
      p10_uge_6774 <= 1'h0;
      p10_uge_6780 <= 1'h0;
      p10_uge_6858 <= 1'h0;
      p10_uge_6938 <= 1'h0;
      p10_uge_7016 <= 1'h0;
      p10_uge_7096 <= 1'h0;
      p10_uge_7102 <= 1'h0;
      p10_uge_7180 <= 1'h0;
      p10_uge_7260 <= 1'h0;
      p10_uge_7338 <= 1'h0;
      p10_r__77 <= 32'h0000_0000;
      p10_bit_slice_6516 <= 1'h0;
      p10_bit_slice_7341 <= 31'h0000_0000;
      p10_bit_slice_6517 <= 1'h0;
      p10_bit_slice_6518 <= 1'h0;
      p10_bit_slice_6519 <= 1'h0;
      p10_bit_slice_6520 <= 1'h0;
      p10_bit_slice_6521 <= 1'h0;
      p10_bit_slice_6522 <= 1'h0;
      p10_bit_slice_6523 <= 1'h0;
      p10_bit_slice_6524 <= 1'h0;
      p10_bit_slice_6525 <= 1'h0;
      p10_bit_slice_6526 <= 1'h0;
      p10_bit_slice_6527 <= 1'h0;
      p10_bit_slice_6528 <= 1'h0;
      p10_bit_slice_6529 <= 1'h0;
      p10_bit_slice_6530 <= 1'h0;
      p10_bit_slice_6531 <= 1'h0;
      p10_bit_slice_6532 <= 1'h0;
      p10_bit_slice_6533 <= 1'h0;
      p10_bit_slice_6534 <= 1'h0;
      p11_b <= 32'h0000_0000;
      p11_uge_6502 <= 1'h0;
      p11_bivisor__1 <= 33'h0_0000_0000;
      p11_uge_6616 <= 1'h0;
      p11_uge_6694 <= 1'h0;
      p11_uge_6774 <= 1'h0;
      p11_uge_6780 <= 1'h0;
      p11_uge_6858 <= 1'h0;
      p11_uge_6938 <= 1'h0;
      p11_uge_7016 <= 1'h0;
      p11_uge_7096 <= 1'h0;
      p11_uge_7102 <= 1'h0;
      p11_uge_7180 <= 1'h0;
      p11_uge_7260 <= 1'h0;
      p11_uge_7338 <= 1'h0;
      p11_uge_7418 <= 1'h0;
      p11_concat_7423 <= 32'h0000_0000;
      p11_uge_7424 <= 1'h0;
      p11_bit_slice_6518 <= 1'h0;
      p11_bit_slice_6519 <= 1'h0;
      p11_bit_slice_6520 <= 1'h0;
      p11_bit_slice_6521 <= 1'h0;
      p11_bit_slice_6522 <= 1'h0;
      p11_bit_slice_6523 <= 1'h0;
      p11_bit_slice_6524 <= 1'h0;
      p11_bit_slice_6525 <= 1'h0;
      p11_bit_slice_6526 <= 1'h0;
      p11_bit_slice_6527 <= 1'h0;
      p11_bit_slice_6528 <= 1'h0;
      p11_bit_slice_6529 <= 1'h0;
      p11_bit_slice_6530 <= 1'h0;
      p11_bit_slice_6531 <= 1'h0;
      p11_bit_slice_6532 <= 1'h0;
      p11_bit_slice_6533 <= 1'h0;
      p11_bit_slice_6534 <= 1'h0;
      p12_b <= 32'h0000_0000;
      p12_uge_6502 <= 1'h0;
      p12_bivisor__1 <= 33'h0_0000_0000;
      p12_uge_6616 <= 1'h0;
      p12_uge_6694 <= 1'h0;
      p12_uge_6774 <= 1'h0;
      p12_uge_6780 <= 1'h0;
      p12_uge_6858 <= 1'h0;
      p12_uge_6938 <= 1'h0;
      p12_uge_7016 <= 1'h0;
      p12_uge_7096 <= 1'h0;
      p12_uge_7102 <= 1'h0;
      p12_uge_7180 <= 1'h0;
      p12_uge_7260 <= 1'h0;
      p12_uge_7338 <= 1'h0;
      p12_uge_7418 <= 1'h0;
      p12_uge_7424 <= 1'h0;
      p12_concat_7501 <= 32'h0000_0000;
      p12_uge_7502 <= 1'h0;
      p12_sub_7503 <= 32'h0000_0000;
      p12_bit_slice_6519 <= 1'h0;
      p12_bit_slice_6520 <= 1'h0;
      p12_bit_slice_6521 <= 1'h0;
      p12_bit_slice_6522 <= 1'h0;
      p12_bit_slice_6523 <= 1'h0;
      p12_bit_slice_6524 <= 1'h0;
      p12_bit_slice_6525 <= 1'h0;
      p12_bit_slice_6526 <= 1'h0;
      p12_bit_slice_6527 <= 1'h0;
      p12_bit_slice_6528 <= 1'h0;
      p12_bit_slice_6529 <= 1'h0;
      p12_bit_slice_6530 <= 1'h0;
      p12_bit_slice_6531 <= 1'h0;
      p12_bit_slice_6532 <= 1'h0;
      p12_bit_slice_6533 <= 1'h0;
      p12_bit_slice_6534 <= 1'h0;
      p13_b <= 32'h0000_0000;
      p13_uge_6502 <= 1'h0;
      p13_bivisor__1 <= 33'h0_0000_0000;
      p13_uge_6616 <= 1'h0;
      p13_uge_6694 <= 1'h0;
      p13_uge_6774 <= 1'h0;
      p13_uge_6780 <= 1'h0;
      p13_uge_6858 <= 1'h0;
      p13_uge_6938 <= 1'h0;
      p13_uge_7016 <= 1'h0;
      p13_uge_7096 <= 1'h0;
      p13_uge_7102 <= 1'h0;
      p13_uge_7180 <= 1'h0;
      p13_uge_7260 <= 1'h0;
      p13_uge_7338 <= 1'h0;
      p13_uge_7418 <= 1'h0;
      p13_uge_7424 <= 1'h0;
      p13_uge_7502 <= 1'h0;
      p13_uge_7582 <= 1'h0;
      p13_r__81 <= 32'h0000_0000;
      p13_bit_slice_6520 <= 1'h0;
      p13_bit_slice_6521 <= 1'h0;
      p13_bit_slice_6522 <= 1'h0;
      p13_bit_slice_6523 <= 1'h0;
      p13_bit_slice_6524 <= 1'h0;
      p13_bit_slice_6525 <= 1'h0;
      p13_bit_slice_6526 <= 1'h0;
      p13_bit_slice_6527 <= 1'h0;
      p13_bit_slice_6528 <= 1'h0;
      p13_bit_slice_6529 <= 1'h0;
      p13_bit_slice_6530 <= 1'h0;
      p13_bit_slice_6531 <= 1'h0;
      p13_bit_slice_6532 <= 1'h0;
      p13_bit_slice_6533 <= 1'h0;
      p13_bit_slice_6534 <= 1'h0;
      p14_b <= 32'h0000_0000;
      p14_uge_6502 <= 1'h0;
      p14_bivisor__1 <= 33'h0_0000_0000;
      p14_uge_6616 <= 1'h0;
      p14_uge_6694 <= 1'h0;
      p14_uge_6774 <= 1'h0;
      p14_uge_6780 <= 1'h0;
      p14_uge_6858 <= 1'h0;
      p14_uge_6938 <= 1'h0;
      p14_uge_7016 <= 1'h0;
      p14_uge_7096 <= 1'h0;
      p14_uge_7102 <= 1'h0;
      p14_uge_7180 <= 1'h0;
      p14_uge_7260 <= 1'h0;
      p14_uge_7338 <= 1'h0;
      p14_uge_7418 <= 1'h0;
      p14_uge_7424 <= 1'h0;
      p14_uge_7502 <= 1'h0;
      p14_uge_7582 <= 1'h0;
      p14_uge_7660 <= 1'h0;
      p14_r__82 <= 32'h0000_0000;
      p14_bit_slice_6521 <= 1'h0;
      p14_bit_slice_7663 <= 31'h0000_0000;
      p14_bit_slice_6522 <= 1'h0;
      p14_bit_slice_6523 <= 1'h0;
      p14_bit_slice_6524 <= 1'h0;
      p14_bit_slice_6525 <= 1'h0;
      p14_bit_slice_6526 <= 1'h0;
      p14_bit_slice_6527 <= 1'h0;
      p14_bit_slice_6528 <= 1'h0;
      p14_bit_slice_6529 <= 1'h0;
      p14_bit_slice_6530 <= 1'h0;
      p14_bit_slice_6531 <= 1'h0;
      p14_bit_slice_6532 <= 1'h0;
      p14_bit_slice_6533 <= 1'h0;
      p14_bit_slice_6534 <= 1'h0;
      p15_b <= 32'h0000_0000;
      p15_uge_6502 <= 1'h0;
      p15_bivisor__1 <= 33'h0_0000_0000;
      p15_uge_6616 <= 1'h0;
      p15_uge_6694 <= 1'h0;
      p15_uge_6774 <= 1'h0;
      p15_uge_6780 <= 1'h0;
      p15_uge_6858 <= 1'h0;
      p15_uge_6938 <= 1'h0;
      p15_uge_7016 <= 1'h0;
      p15_uge_7096 <= 1'h0;
      p15_uge_7102 <= 1'h0;
      p15_uge_7180 <= 1'h0;
      p15_uge_7260 <= 1'h0;
      p15_uge_7338 <= 1'h0;
      p15_uge_7418 <= 1'h0;
      p15_uge_7424 <= 1'h0;
      p15_uge_7502 <= 1'h0;
      p15_uge_7582 <= 1'h0;
      p15_uge_7660 <= 1'h0;
      p15_uge_7740 <= 1'h0;
      p15_concat_7745 <= 32'h0000_0000;
      p15_uge_7746 <= 1'h0;
      p15_bit_slice_6523 <= 1'h0;
      p15_bit_slice_6524 <= 1'h0;
      p15_bit_slice_6525 <= 1'h0;
      p15_bit_slice_6526 <= 1'h0;
      p15_bit_slice_6527 <= 1'h0;
      p15_bit_slice_6528 <= 1'h0;
      p15_bit_slice_6529 <= 1'h0;
      p15_bit_slice_6530 <= 1'h0;
      p15_bit_slice_6531 <= 1'h0;
      p15_bit_slice_6532 <= 1'h0;
      p15_bit_slice_6533 <= 1'h0;
      p15_bit_slice_6534 <= 1'h0;
      p16_b <= 32'h0000_0000;
      p16_uge_6502 <= 1'h0;
      p16_bivisor__1 <= 33'h0_0000_0000;
      p16_uge_6616 <= 1'h0;
      p16_uge_6694 <= 1'h0;
      p16_uge_6774 <= 1'h0;
      p16_uge_6780 <= 1'h0;
      p16_uge_6858 <= 1'h0;
      p16_uge_6938 <= 1'h0;
      p16_uge_7016 <= 1'h0;
      p16_uge_7096 <= 1'h0;
      p16_uge_7102 <= 1'h0;
      p16_uge_7180 <= 1'h0;
      p16_uge_7260 <= 1'h0;
      p16_uge_7338 <= 1'h0;
      p16_uge_7418 <= 1'h0;
      p16_uge_7424 <= 1'h0;
      p16_uge_7502 <= 1'h0;
      p16_uge_7582 <= 1'h0;
      p16_uge_7660 <= 1'h0;
      p16_uge_7740 <= 1'h0;
      p16_uge_7746 <= 1'h0;
      p16_concat_7823 <= 32'h0000_0000;
      p16_uge_7824 <= 1'h0;
      p16_sub_7825 <= 32'h0000_0000;
      p16_bit_slice_6524 <= 1'h0;
      p16_bit_slice_6525 <= 1'h0;
      p16_bit_slice_6526 <= 1'h0;
      p16_bit_slice_6527 <= 1'h0;
      p16_bit_slice_6528 <= 1'h0;
      p16_bit_slice_6529 <= 1'h0;
      p16_bit_slice_6530 <= 1'h0;
      p16_bit_slice_6531 <= 1'h0;
      p16_bit_slice_6532 <= 1'h0;
      p16_bit_slice_6533 <= 1'h0;
      p16_bit_slice_6534 <= 1'h0;
      p17_b <= 32'h0000_0000;
      p17_uge_6502 <= 1'h0;
      p17_bivisor__1 <= 33'h0_0000_0000;
      p17_uge_6616 <= 1'h0;
      p17_uge_6694 <= 1'h0;
      p17_uge_6774 <= 1'h0;
      p17_uge_6780 <= 1'h0;
      p17_uge_6858 <= 1'h0;
      p17_uge_6938 <= 1'h0;
      p17_uge_7016 <= 1'h0;
      p17_uge_7096 <= 1'h0;
      p17_uge_7102 <= 1'h0;
      p17_uge_7180 <= 1'h0;
      p17_uge_7260 <= 1'h0;
      p17_uge_7338 <= 1'h0;
      p17_uge_7418 <= 1'h0;
      p17_uge_7424 <= 1'h0;
      p17_uge_7502 <= 1'h0;
      p17_uge_7582 <= 1'h0;
      p17_uge_7660 <= 1'h0;
      p17_uge_7740 <= 1'h0;
      p17_uge_7746 <= 1'h0;
      p17_uge_7824 <= 1'h0;
      p17_uge_7904 <= 1'h0;
      p17_r__86 <= 32'h0000_0000;
      p17_bit_slice_6525 <= 1'h0;
      p17_bit_slice_6526 <= 1'h0;
      p17_bit_slice_6527 <= 1'h0;
      p17_bit_slice_6528 <= 1'h0;
      p17_bit_slice_6529 <= 1'h0;
      p17_bit_slice_6530 <= 1'h0;
      p17_bit_slice_6531 <= 1'h0;
      p17_bit_slice_6532 <= 1'h0;
      p17_bit_slice_6533 <= 1'h0;
      p17_bit_slice_6534 <= 1'h0;
      p18_b <= 32'h0000_0000;
      p18_uge_6502 <= 1'h0;
      p18_bivisor__1 <= 33'h0_0000_0000;
      p18_uge_6616 <= 1'h0;
      p18_uge_6694 <= 1'h0;
      p18_uge_6774 <= 1'h0;
      p18_uge_6780 <= 1'h0;
      p18_uge_6858 <= 1'h0;
      p18_uge_6938 <= 1'h0;
      p18_uge_7016 <= 1'h0;
      p18_uge_7096 <= 1'h0;
      p18_uge_7102 <= 1'h0;
      p18_uge_7180 <= 1'h0;
      p18_uge_7260 <= 1'h0;
      p18_uge_7338 <= 1'h0;
      p18_uge_7418 <= 1'h0;
      p18_uge_7424 <= 1'h0;
      p18_uge_7502 <= 1'h0;
      p18_uge_7582 <= 1'h0;
      p18_uge_7660 <= 1'h0;
      p18_uge_7740 <= 1'h0;
      p18_uge_7746 <= 1'h0;
      p18_uge_7824 <= 1'h0;
      p18_uge_7904 <= 1'h0;
      p18_uge_7982 <= 1'h0;
      p18_r__87 <= 32'h0000_0000;
      p18_bit_slice_6526 <= 1'h0;
      p18_bit_slice_7985 <= 31'h0000_0000;
      p18_bit_slice_6527 <= 1'h0;
      p18_bit_slice_6528 <= 1'h0;
      p18_bit_slice_6529 <= 1'h0;
      p18_bit_slice_6530 <= 1'h0;
      p18_bit_slice_6531 <= 1'h0;
      p18_bit_slice_6532 <= 1'h0;
      p18_bit_slice_6533 <= 1'h0;
      p18_bit_slice_6534 <= 1'h0;
      p19_b <= 32'h0000_0000;
      p19_uge_6502 <= 1'h0;
      p19_bivisor__1 <= 33'h0_0000_0000;
      p19_uge_6616 <= 1'h0;
      p19_uge_6694 <= 1'h0;
      p19_uge_6774 <= 1'h0;
      p19_uge_6780 <= 1'h0;
      p19_uge_6858 <= 1'h0;
      p19_uge_6938 <= 1'h0;
      p19_uge_7016 <= 1'h0;
      p19_uge_7096 <= 1'h0;
      p19_uge_7102 <= 1'h0;
      p19_uge_7180 <= 1'h0;
      p19_uge_7260 <= 1'h0;
      p19_uge_7338 <= 1'h0;
      p19_uge_7418 <= 1'h0;
      p19_uge_7424 <= 1'h0;
      p19_uge_7502 <= 1'h0;
      p19_uge_7582 <= 1'h0;
      p19_uge_7660 <= 1'h0;
      p19_uge_7740 <= 1'h0;
      p19_uge_7746 <= 1'h0;
      p19_uge_7824 <= 1'h0;
      p19_uge_7904 <= 1'h0;
      p19_uge_7982 <= 1'h0;
      p19_uge_8062 <= 1'h0;
      p19_concat_8067 <= 32'h0000_0000;
      p19_uge_8068 <= 1'h0;
      p19_bit_slice_6528 <= 1'h0;
      p19_bit_slice_6529 <= 1'h0;
      p19_bit_slice_6530 <= 1'h0;
      p19_bit_slice_6531 <= 1'h0;
      p19_bit_slice_6532 <= 1'h0;
      p19_bit_slice_6533 <= 1'h0;
      p19_bit_slice_6534 <= 1'h0;
      p20_b <= 32'h0000_0000;
      p20_uge_6502 <= 1'h0;
      p20_bivisor__1 <= 33'h0_0000_0000;
      p20_uge_6616 <= 1'h0;
      p20_uge_6694 <= 1'h0;
      p20_uge_6774 <= 1'h0;
      p20_uge_6780 <= 1'h0;
      p20_uge_6858 <= 1'h0;
      p20_uge_6938 <= 1'h0;
      p20_uge_7016 <= 1'h0;
      p20_uge_7096 <= 1'h0;
      p20_uge_7102 <= 1'h0;
      p20_uge_7180 <= 1'h0;
      p20_uge_7260 <= 1'h0;
      p20_uge_7338 <= 1'h0;
      p20_uge_7418 <= 1'h0;
      p20_uge_7424 <= 1'h0;
      p20_uge_7502 <= 1'h0;
      p20_uge_7582 <= 1'h0;
      p20_uge_7660 <= 1'h0;
      p20_uge_7740 <= 1'h0;
      p20_uge_7746 <= 1'h0;
      p20_uge_7824 <= 1'h0;
      p20_uge_7904 <= 1'h0;
      p20_uge_7982 <= 1'h0;
      p20_uge_8062 <= 1'h0;
      p20_uge_8068 <= 1'h0;
      p20_concat_8145 <= 32'h0000_0000;
      p20_uge_8146 <= 1'h0;
      p20_sub_8147 <= 32'h0000_0000;
      p20_bit_slice_6529 <= 1'h0;
      p20_bit_slice_6530 <= 1'h0;
      p20_bit_slice_6531 <= 1'h0;
      p20_bit_slice_6532 <= 1'h0;
      p20_bit_slice_6533 <= 1'h0;
      p20_bit_slice_6534 <= 1'h0;
      p21_b <= 32'h0000_0000;
      p21_uge_6502 <= 1'h0;
      p21_bivisor__1 <= 33'h0_0000_0000;
      p21_uge_6616 <= 1'h0;
      p21_uge_6694 <= 1'h0;
      p21_uge_6774 <= 1'h0;
      p21_uge_6780 <= 1'h0;
      p21_uge_6858 <= 1'h0;
      p21_uge_6938 <= 1'h0;
      p21_uge_7016 <= 1'h0;
      p21_uge_7096 <= 1'h0;
      p21_uge_7102 <= 1'h0;
      p21_uge_7180 <= 1'h0;
      p21_uge_7260 <= 1'h0;
      p21_uge_7338 <= 1'h0;
      p21_uge_7418 <= 1'h0;
      p21_uge_7424 <= 1'h0;
      p21_uge_7502 <= 1'h0;
      p21_uge_7582 <= 1'h0;
      p21_uge_7660 <= 1'h0;
      p21_uge_7740 <= 1'h0;
      p21_uge_7746 <= 1'h0;
      p21_uge_7824 <= 1'h0;
      p21_uge_7904 <= 1'h0;
      p21_uge_7982 <= 1'h0;
      p21_uge_8062 <= 1'h0;
      p21_uge_8068 <= 1'h0;
      p21_uge_8146 <= 1'h0;
      p21_uge_8226 <= 1'h0;
      p21_r__91 <= 32'h0000_0000;
      p21_bit_slice_6530 <= 1'h0;
      p21_bit_slice_6531 <= 1'h0;
      p21_bit_slice_6532 <= 1'h0;
      p21_bit_slice_6533 <= 1'h0;
      p21_bit_slice_6534 <= 1'h0;
      p22_b <= 32'h0000_0000;
      p22_uge_6502 <= 1'h0;
      p22_bivisor__1 <= 33'h0_0000_0000;
      p22_uge_6616 <= 1'h0;
      p22_uge_6694 <= 1'h0;
      p22_uge_6774 <= 1'h0;
      p22_uge_6780 <= 1'h0;
      p22_uge_6858 <= 1'h0;
      p22_uge_6938 <= 1'h0;
      p22_uge_7016 <= 1'h0;
      p22_uge_7096 <= 1'h0;
      p22_uge_7102 <= 1'h0;
      p22_uge_7180 <= 1'h0;
      p22_uge_7260 <= 1'h0;
      p22_uge_7338 <= 1'h0;
      p22_uge_7418 <= 1'h0;
      p22_uge_7424 <= 1'h0;
      p22_uge_7502 <= 1'h0;
      p22_uge_7582 <= 1'h0;
      p22_uge_7660 <= 1'h0;
      p22_uge_7740 <= 1'h0;
      p22_uge_7746 <= 1'h0;
      p22_uge_7824 <= 1'h0;
      p22_uge_7904 <= 1'h0;
      p22_uge_7982 <= 1'h0;
      p22_uge_8062 <= 1'h0;
      p22_uge_8068 <= 1'h0;
      p22_uge_8146 <= 1'h0;
      p22_uge_8226 <= 1'h0;
      p22_uge_8304 <= 1'h0;
      p22_r__92 <= 32'h0000_0000;
      p22_bit_slice_6531 <= 1'h0;
      p22_bit_slice_8307 <= 31'h0000_0000;
      p22_bit_slice_6532 <= 1'h0;
      p22_bit_slice_6533 <= 1'h0;
      p22_bit_slice_6534 <= 1'h0;
      p23_b <= 32'h0000_0000;
      p23_uge_6502 <= 1'h0;
      p23_bivisor__1 <= 33'h0_0000_0000;
      p23_uge_6616 <= 1'h0;
      p23_uge_6694 <= 1'h0;
      p23_uge_6774 <= 1'h0;
      p23_uge_6780 <= 1'h0;
      p23_uge_6858 <= 1'h0;
      p23_uge_6938 <= 1'h0;
      p23_uge_7016 <= 1'h0;
      p23_uge_7096 <= 1'h0;
      p23_uge_7102 <= 1'h0;
      p23_uge_7180 <= 1'h0;
      p23_uge_7260 <= 1'h0;
      p23_uge_7338 <= 1'h0;
      p23_uge_7418 <= 1'h0;
      p23_uge_7424 <= 1'h0;
      p23_uge_7502 <= 1'h0;
      p23_uge_7582 <= 1'h0;
      p23_uge_7660 <= 1'h0;
      p23_uge_7740 <= 1'h0;
      p23_uge_7746 <= 1'h0;
      p23_uge_7824 <= 1'h0;
      p23_uge_7904 <= 1'h0;
      p23_uge_7982 <= 1'h0;
      p23_uge_8062 <= 1'h0;
      p23_uge_8068 <= 1'h0;
      p23_uge_8146 <= 1'h0;
      p23_uge_8226 <= 1'h0;
      p23_uge_8304 <= 1'h0;
      p23_uge_8384 <= 1'h0;
      p23_concat_8389 <= 32'h0000_0000;
      p23_uge_8390 <= 1'h0;
      p23_bit_slice_6533 <= 1'h0;
      p23_bit_slice_6534 <= 1'h0;
      p24_uge_6502 <= 1'h0;
      p24_bivisor__1 <= 33'h0_0000_0000;
      p24_uge_6616 <= 1'h0;
      p24_uge_6694 <= 1'h0;
      p24_uge_6774 <= 1'h0;
      p24_uge_6780 <= 1'h0;
      p24_uge_6858 <= 1'h0;
      p24_uge_6938 <= 1'h0;
      p24_uge_7016 <= 1'h0;
      p24_uge_7096 <= 1'h0;
      p24_uge_7102 <= 1'h0;
      p24_uge_7180 <= 1'h0;
      p24_uge_7260 <= 1'h0;
      p24_uge_7338 <= 1'h0;
      p24_uge_7418 <= 1'h0;
      p24_uge_7424 <= 1'h0;
      p24_uge_7502 <= 1'h0;
      p24_uge_7582 <= 1'h0;
      p24_uge_7660 <= 1'h0;
      p24_uge_7740 <= 1'h0;
      p24_uge_7746 <= 1'h0;
      p24_uge_7824 <= 1'h0;
      p24_uge_7904 <= 1'h0;
      p24_uge_7982 <= 1'h0;
      p24_uge_8062 <= 1'h0;
      p24_uge_8068 <= 1'h0;
      p24_uge_8146 <= 1'h0;
      p24_uge_8226 <= 1'h0;
      p24_uge_8304 <= 1'h0;
      p24_uge_8384 <= 1'h0;
      p24_uge_8390 <= 1'h0;
      p24_concat_8467 <= 32'h0000_0000;
      p24_uge_8468 <= 1'h0;
      p24_sub_8469 <= 32'h0000_0000;
      p24_bit_slice_6534 <= 1'h0;
      p0_valid <= 1'h0;
      p1_valid <= 1'h0;
      p2_valid <= 1'h0;
      p3_valid <= 1'h0;
      p4_valid <= 1'h0;
      p5_valid <= 1'h0;
      p6_valid <= 1'h0;
      p7_valid <= 1'h0;
      p8_valid <= 1'h0;
      p9_valid <= 1'h0;
      p10_valid <= 1'h0;
      p11_valid <= 1'h0;
      p12_valid <= 1'h0;
      p13_valid <= 1'h0;
      p14_valid <= 1'h0;
      p15_valid <= 1'h0;
      p16_valid <= 1'h0;
      p17_valid <= 1'h0;
      p18_valid <= 1'h0;
      p19_valid <= 1'h0;
      p20_valid <= 1'h0;
      p21_valid <= 1'h0;
      p22_valid <= 1'h0;
      p23_valid <= 1'h0;
      p24_valid <= 1'h0;
      p25_valid <= 1'h0;
      p26_valid <= 1'h0;
      p27_valid <= 1'h0;
      p28_valid <= 1'h0;
      p29_valid <= 1'h0;
      p30_valid <= 1'h0;
      lhs_reg <= 32'h0000_0000;
      lhs_valid_reg <= 1'h0;
      rhs_reg <= 32'h0000_0000;
      rhs_valid_reg <= 1'h0;
      result_reg <= 32'h0000_0000;
      result_valid_reg <= 1'h0;
    end else begin
      p0_concat_6500 <= p0_data_enable ? concat_6500 : p0_concat_6500;
      p0_b <= p0_data_enable ? rhs_reg : p0_b;
      p0_uge_6502 <= p0_data_enable ? uge_6502 : p0_uge_6502;
      p0_sub_6503 <= p0_data_enable ? sub_6503 : p0_sub_6503;
      p0_bit_slice_6504 <= p0_data_enable ? bit_slice_6504 : p0_bit_slice_6504;
      p0_bit_slice_6505 <= p0_data_enable ? bit_slice_6505 : p0_bit_slice_6505;
      p0_bit_slice_6506 <= p0_data_enable ? bit_slice_6506 : p0_bit_slice_6506;
      p0_bit_slice_6507 <= p0_data_enable ? bit_slice_6507 : p0_bit_slice_6507;
      p0_bit_slice_6508 <= p0_data_enable ? bit_slice_6508 : p0_bit_slice_6508;
      p0_bit_slice_6509 <= p0_data_enable ? bit_slice_6509 : p0_bit_slice_6509;
      p0_bit_slice_6510 <= p0_data_enable ? bit_slice_6510 : p0_bit_slice_6510;
      p0_bit_slice_6511 <= p0_data_enable ? bit_slice_6511 : p0_bit_slice_6511;
      p0_bit_slice_6512 <= p0_data_enable ? bit_slice_6512 : p0_bit_slice_6512;
      p0_bit_slice_6513 <= p0_data_enable ? bit_slice_6513 : p0_bit_slice_6513;
      p0_bit_slice_6514 <= p0_data_enable ? bit_slice_6514 : p0_bit_slice_6514;
      p0_bit_slice_6515 <= p0_data_enable ? bit_slice_6515 : p0_bit_slice_6515;
      p0_bit_slice_6516 <= p0_data_enable ? bit_slice_6516 : p0_bit_slice_6516;
      p0_bit_slice_6517 <= p0_data_enable ? bit_slice_6517 : p0_bit_slice_6517;
      p0_bit_slice_6518 <= p0_data_enable ? bit_slice_6518 : p0_bit_slice_6518;
      p0_bit_slice_6519 <= p0_data_enable ? bit_slice_6519 : p0_bit_slice_6519;
      p0_bit_slice_6520 <= p0_data_enable ? bit_slice_6520 : p0_bit_slice_6520;
      p0_bit_slice_6521 <= p0_data_enable ? bit_slice_6521 : p0_bit_slice_6521;
      p0_bit_slice_6522 <= p0_data_enable ? bit_slice_6522 : p0_bit_slice_6522;
      p0_bit_slice_6523 <= p0_data_enable ? bit_slice_6523 : p0_bit_slice_6523;
      p0_bit_slice_6524 <= p0_data_enable ? bit_slice_6524 : p0_bit_slice_6524;
      p0_bit_slice_6525 <= p0_data_enable ? bit_slice_6525 : p0_bit_slice_6525;
      p0_bit_slice_6526 <= p0_data_enable ? bit_slice_6526 : p0_bit_slice_6526;
      p0_bit_slice_6527 <= p0_data_enable ? bit_slice_6527 : p0_bit_slice_6527;
      p0_bit_slice_6528 <= p0_data_enable ? bit_slice_6528 : p0_bit_slice_6528;
      p0_bit_slice_6529 <= p0_data_enable ? bit_slice_6529 : p0_bit_slice_6529;
      p0_bit_slice_6530 <= p0_data_enable ? bit_slice_6530 : p0_bit_slice_6530;
      p0_bit_slice_6531 <= p0_data_enable ? bit_slice_6531 : p0_bit_slice_6531;
      p0_bit_slice_6532 <= p0_data_enable ? bit_slice_6532 : p0_bit_slice_6532;
      p0_bit_slice_6533 <= p0_data_enable ? bit_slice_6533 : p0_bit_slice_6533;
      p0_bit_slice_6534 <= p0_data_enable ? bit_slice_6534 : p0_bit_slice_6534;
      p1_b <= p1_data_enable ? p0_b : p1_b;
      p1_uge_6502 <= p1_data_enable ? p0_uge_6502 : p1_uge_6502;
      p1_bivisor__1 <= p1_data_enable ? bivisor__1 : p1_bivisor__1;
      p1_uge_6616 <= p1_data_enable ? uge_6616 : p1_uge_6616;
      p1_r__66 <= p1_data_enable ? r__66 : p1_r__66;
      p1_bit_slice_6505 <= p1_data_enable ? p0_bit_slice_6505 : p1_bit_slice_6505;
      p1_bit_slice_6506 <= p1_data_enable ? p0_bit_slice_6506 : p1_bit_slice_6506;
      p1_bit_slice_6507 <= p1_data_enable ? p0_bit_slice_6507 : p1_bit_slice_6507;
      p1_bit_slice_6508 <= p1_data_enable ? p0_bit_slice_6508 : p1_bit_slice_6508;
      p1_bit_slice_6509 <= p1_data_enable ? p0_bit_slice_6509 : p1_bit_slice_6509;
      p1_bit_slice_6510 <= p1_data_enable ? p0_bit_slice_6510 : p1_bit_slice_6510;
      p1_bit_slice_6511 <= p1_data_enable ? p0_bit_slice_6511 : p1_bit_slice_6511;
      p1_bit_slice_6512 <= p1_data_enable ? p0_bit_slice_6512 : p1_bit_slice_6512;
      p1_bit_slice_6513 <= p1_data_enable ? p0_bit_slice_6513 : p1_bit_slice_6513;
      p1_bit_slice_6514 <= p1_data_enable ? p0_bit_slice_6514 : p1_bit_slice_6514;
      p1_bit_slice_6515 <= p1_data_enable ? p0_bit_slice_6515 : p1_bit_slice_6515;
      p1_bit_slice_6516 <= p1_data_enable ? p0_bit_slice_6516 : p1_bit_slice_6516;
      p1_bit_slice_6517 <= p1_data_enable ? p0_bit_slice_6517 : p1_bit_slice_6517;
      p1_bit_slice_6518 <= p1_data_enable ? p0_bit_slice_6518 : p1_bit_slice_6518;
      p1_bit_slice_6519 <= p1_data_enable ? p0_bit_slice_6519 : p1_bit_slice_6519;
      p1_bit_slice_6520 <= p1_data_enable ? p0_bit_slice_6520 : p1_bit_slice_6520;
      p1_bit_slice_6521 <= p1_data_enable ? p0_bit_slice_6521 : p1_bit_slice_6521;
      p1_bit_slice_6522 <= p1_data_enable ? p0_bit_slice_6522 : p1_bit_slice_6522;
      p1_bit_slice_6523 <= p1_data_enable ? p0_bit_slice_6523 : p1_bit_slice_6523;
      p1_bit_slice_6524 <= p1_data_enable ? p0_bit_slice_6524 : p1_bit_slice_6524;
      p1_bit_slice_6525 <= p1_data_enable ? p0_bit_slice_6525 : p1_bit_slice_6525;
      p1_bit_slice_6526 <= p1_data_enable ? p0_bit_slice_6526 : p1_bit_slice_6526;
      p1_bit_slice_6527 <= p1_data_enable ? p0_bit_slice_6527 : p1_bit_slice_6527;
      p1_bit_slice_6528 <= p1_data_enable ? p0_bit_slice_6528 : p1_bit_slice_6528;
      p1_bit_slice_6529 <= p1_data_enable ? p0_bit_slice_6529 : p1_bit_slice_6529;
      p1_bit_slice_6530 <= p1_data_enable ? p0_bit_slice_6530 : p1_bit_slice_6530;
      p1_bit_slice_6531 <= p1_data_enable ? p0_bit_slice_6531 : p1_bit_slice_6531;
      p1_bit_slice_6532 <= p1_data_enable ? p0_bit_slice_6532 : p1_bit_slice_6532;
      p1_bit_slice_6533 <= p1_data_enable ? p0_bit_slice_6533 : p1_bit_slice_6533;
      p1_bit_slice_6534 <= p1_data_enable ? p0_bit_slice_6534 : p1_bit_slice_6534;
      p2_b <= p2_data_enable ? p1_b : p2_b;
      p2_uge_6502 <= p2_data_enable ? p1_uge_6502 : p2_uge_6502;
      p2_bivisor__1 <= p2_data_enable ? p1_bivisor__1 : p2_bivisor__1;
      p2_uge_6616 <= p2_data_enable ? p1_uge_6616 : p2_uge_6616;
      p2_uge_6694 <= p2_data_enable ? uge_6694 : p2_uge_6694;
      p2_r__67 <= p2_data_enable ? r__67 : p2_r__67;
      p2_bit_slice_6506 <= p2_data_enable ? p1_bit_slice_6506 : p2_bit_slice_6506;
      p2_bit_slice_6697 <= p2_data_enable ? bit_slice_6697 : p2_bit_slice_6697;
      p2_bit_slice_6507 <= p2_data_enable ? p1_bit_slice_6507 : p2_bit_slice_6507;
      p2_bit_slice_6508 <= p2_data_enable ? p1_bit_slice_6508 : p2_bit_slice_6508;
      p2_bit_slice_6509 <= p2_data_enable ? p1_bit_slice_6509 : p2_bit_slice_6509;
      p2_bit_slice_6510 <= p2_data_enable ? p1_bit_slice_6510 : p2_bit_slice_6510;
      p2_bit_slice_6511 <= p2_data_enable ? p1_bit_slice_6511 : p2_bit_slice_6511;
      p2_bit_slice_6512 <= p2_data_enable ? p1_bit_slice_6512 : p2_bit_slice_6512;
      p2_bit_slice_6513 <= p2_data_enable ? p1_bit_slice_6513 : p2_bit_slice_6513;
      p2_bit_slice_6514 <= p2_data_enable ? p1_bit_slice_6514 : p2_bit_slice_6514;
      p2_bit_slice_6515 <= p2_data_enable ? p1_bit_slice_6515 : p2_bit_slice_6515;
      p2_bit_slice_6516 <= p2_data_enable ? p1_bit_slice_6516 : p2_bit_slice_6516;
      p2_bit_slice_6517 <= p2_data_enable ? p1_bit_slice_6517 : p2_bit_slice_6517;
      p2_bit_slice_6518 <= p2_data_enable ? p1_bit_slice_6518 : p2_bit_slice_6518;
      p2_bit_slice_6519 <= p2_data_enable ? p1_bit_slice_6519 : p2_bit_slice_6519;
      p2_bit_slice_6520 <= p2_data_enable ? p1_bit_slice_6520 : p2_bit_slice_6520;
      p2_bit_slice_6521 <= p2_data_enable ? p1_bit_slice_6521 : p2_bit_slice_6521;
      p2_bit_slice_6522 <= p2_data_enable ? p1_bit_slice_6522 : p2_bit_slice_6522;
      p2_bit_slice_6523 <= p2_data_enable ? p1_bit_slice_6523 : p2_bit_slice_6523;
      p2_bit_slice_6524 <= p2_data_enable ? p1_bit_slice_6524 : p2_bit_slice_6524;
      p2_bit_slice_6525 <= p2_data_enable ? p1_bit_slice_6525 : p2_bit_slice_6525;
      p2_bit_slice_6526 <= p2_data_enable ? p1_bit_slice_6526 : p2_bit_slice_6526;
      p2_bit_slice_6527 <= p2_data_enable ? p1_bit_slice_6527 : p2_bit_slice_6527;
      p2_bit_slice_6528 <= p2_data_enable ? p1_bit_slice_6528 : p2_bit_slice_6528;
      p2_bit_slice_6529 <= p2_data_enable ? p1_bit_slice_6529 : p2_bit_slice_6529;
      p2_bit_slice_6530 <= p2_data_enable ? p1_bit_slice_6530 : p2_bit_slice_6530;
      p2_bit_slice_6531 <= p2_data_enable ? p1_bit_slice_6531 : p2_bit_slice_6531;
      p2_bit_slice_6532 <= p2_data_enable ? p1_bit_slice_6532 : p2_bit_slice_6532;
      p2_bit_slice_6533 <= p2_data_enable ? p1_bit_slice_6533 : p2_bit_slice_6533;
      p2_bit_slice_6534 <= p2_data_enable ? p1_bit_slice_6534 : p2_bit_slice_6534;
      p3_b <= p3_data_enable ? p2_b : p3_b;
      p3_uge_6502 <= p3_data_enable ? p2_uge_6502 : p3_uge_6502;
      p3_bivisor__1 <= p3_data_enable ? p2_bivisor__1 : p3_bivisor__1;
      p3_uge_6616 <= p3_data_enable ? p2_uge_6616 : p3_uge_6616;
      p3_uge_6694 <= p3_data_enable ? p2_uge_6694 : p3_uge_6694;
      p3_uge_6774 <= p3_data_enable ? uge_6774 : p3_uge_6774;
      p3_concat_6779 <= p3_data_enable ? concat_6779 : p3_concat_6779;
      p3_uge_6780 <= p3_data_enable ? uge_6780 : p3_uge_6780;
      p3_bit_slice_6508 <= p3_data_enable ? p2_bit_slice_6508 : p3_bit_slice_6508;
      p3_bit_slice_6509 <= p3_data_enable ? p2_bit_slice_6509 : p3_bit_slice_6509;
      p3_bit_slice_6510 <= p3_data_enable ? p2_bit_slice_6510 : p3_bit_slice_6510;
      p3_bit_slice_6511 <= p3_data_enable ? p2_bit_slice_6511 : p3_bit_slice_6511;
      p3_bit_slice_6512 <= p3_data_enable ? p2_bit_slice_6512 : p3_bit_slice_6512;
      p3_bit_slice_6513 <= p3_data_enable ? p2_bit_slice_6513 : p3_bit_slice_6513;
      p3_bit_slice_6514 <= p3_data_enable ? p2_bit_slice_6514 : p3_bit_slice_6514;
      p3_bit_slice_6515 <= p3_data_enable ? p2_bit_slice_6515 : p3_bit_slice_6515;
      p3_bit_slice_6516 <= p3_data_enable ? p2_bit_slice_6516 : p3_bit_slice_6516;
      p3_bit_slice_6517 <= p3_data_enable ? p2_bit_slice_6517 : p3_bit_slice_6517;
      p3_bit_slice_6518 <= p3_data_enable ? p2_bit_slice_6518 : p3_bit_slice_6518;
      p3_bit_slice_6519 <= p3_data_enable ? p2_bit_slice_6519 : p3_bit_slice_6519;
      p3_bit_slice_6520 <= p3_data_enable ? p2_bit_slice_6520 : p3_bit_slice_6520;
      p3_bit_slice_6521 <= p3_data_enable ? p2_bit_slice_6521 : p3_bit_slice_6521;
      p3_bit_slice_6522 <= p3_data_enable ? p2_bit_slice_6522 : p3_bit_slice_6522;
      p3_bit_slice_6523 <= p3_data_enable ? p2_bit_slice_6523 : p3_bit_slice_6523;
      p3_bit_slice_6524 <= p3_data_enable ? p2_bit_slice_6524 : p3_bit_slice_6524;
      p3_bit_slice_6525 <= p3_data_enable ? p2_bit_slice_6525 : p3_bit_slice_6525;
      p3_bit_slice_6526 <= p3_data_enable ? p2_bit_slice_6526 : p3_bit_slice_6526;
      p3_bit_slice_6527 <= p3_data_enable ? p2_bit_slice_6527 : p3_bit_slice_6527;
      p3_bit_slice_6528 <= p3_data_enable ? p2_bit_slice_6528 : p3_bit_slice_6528;
      p3_bit_slice_6529 <= p3_data_enable ? p2_bit_slice_6529 : p3_bit_slice_6529;
      p3_bit_slice_6530 <= p3_data_enable ? p2_bit_slice_6530 : p3_bit_slice_6530;
      p3_bit_slice_6531 <= p3_data_enable ? p2_bit_slice_6531 : p3_bit_slice_6531;
      p3_bit_slice_6532 <= p3_data_enable ? p2_bit_slice_6532 : p3_bit_slice_6532;
      p3_bit_slice_6533 <= p3_data_enable ? p2_bit_slice_6533 : p3_bit_slice_6533;
      p3_bit_slice_6534 <= p3_data_enable ? p2_bit_slice_6534 : p3_bit_slice_6534;
      p4_b <= p4_data_enable ? p3_b : p4_b;
      p4_uge_6502 <= p4_data_enable ? p3_uge_6502 : p4_uge_6502;
      p4_bivisor__1 <= p4_data_enable ? p3_bivisor__1 : p4_bivisor__1;
      p4_uge_6616 <= p4_data_enable ? p3_uge_6616 : p4_uge_6616;
      p4_uge_6694 <= p4_data_enable ? p3_uge_6694 : p4_uge_6694;
      p4_uge_6774 <= p4_data_enable ? p3_uge_6774 : p4_uge_6774;
      p4_uge_6780 <= p4_data_enable ? p3_uge_6780 : p4_uge_6780;
      p4_concat_6857 <= p4_data_enable ? concat_6857 : p4_concat_6857;
      p4_uge_6858 <= p4_data_enable ? uge_6858 : p4_uge_6858;
      p4_sub_6859 <= p4_data_enable ? sub_6859 : p4_sub_6859;
      p4_bit_slice_6509 <= p4_data_enable ? p3_bit_slice_6509 : p4_bit_slice_6509;
      p4_bit_slice_6510 <= p4_data_enable ? p3_bit_slice_6510 : p4_bit_slice_6510;
      p4_bit_slice_6511 <= p4_data_enable ? p3_bit_slice_6511 : p4_bit_slice_6511;
      p4_bit_slice_6512 <= p4_data_enable ? p3_bit_slice_6512 : p4_bit_slice_6512;
      p4_bit_slice_6513 <= p4_data_enable ? p3_bit_slice_6513 : p4_bit_slice_6513;
      p4_bit_slice_6514 <= p4_data_enable ? p3_bit_slice_6514 : p4_bit_slice_6514;
      p4_bit_slice_6515 <= p4_data_enable ? p3_bit_slice_6515 : p4_bit_slice_6515;
      p4_bit_slice_6516 <= p4_data_enable ? p3_bit_slice_6516 : p4_bit_slice_6516;
      p4_bit_slice_6517 <= p4_data_enable ? p3_bit_slice_6517 : p4_bit_slice_6517;
      p4_bit_slice_6518 <= p4_data_enable ? p3_bit_slice_6518 : p4_bit_slice_6518;
      p4_bit_slice_6519 <= p4_data_enable ? p3_bit_slice_6519 : p4_bit_slice_6519;
      p4_bit_slice_6520 <= p4_data_enable ? p3_bit_slice_6520 : p4_bit_slice_6520;
      p4_bit_slice_6521 <= p4_data_enable ? p3_bit_slice_6521 : p4_bit_slice_6521;
      p4_bit_slice_6522 <= p4_data_enable ? p3_bit_slice_6522 : p4_bit_slice_6522;
      p4_bit_slice_6523 <= p4_data_enable ? p3_bit_slice_6523 : p4_bit_slice_6523;
      p4_bit_slice_6524 <= p4_data_enable ? p3_bit_slice_6524 : p4_bit_slice_6524;
      p4_bit_slice_6525 <= p4_data_enable ? p3_bit_slice_6525 : p4_bit_slice_6525;
      p4_bit_slice_6526 <= p4_data_enable ? p3_bit_slice_6526 : p4_bit_slice_6526;
      p4_bit_slice_6527 <= p4_data_enable ? p3_bit_slice_6527 : p4_bit_slice_6527;
      p4_bit_slice_6528 <= p4_data_enable ? p3_bit_slice_6528 : p4_bit_slice_6528;
      p4_bit_slice_6529 <= p4_data_enable ? p3_bit_slice_6529 : p4_bit_slice_6529;
      p4_bit_slice_6530 <= p4_data_enable ? p3_bit_slice_6530 : p4_bit_slice_6530;
      p4_bit_slice_6531 <= p4_data_enable ? p3_bit_slice_6531 : p4_bit_slice_6531;
      p4_bit_slice_6532 <= p4_data_enable ? p3_bit_slice_6532 : p4_bit_slice_6532;
      p4_bit_slice_6533 <= p4_data_enable ? p3_bit_slice_6533 : p4_bit_slice_6533;
      p4_bit_slice_6534 <= p4_data_enable ? p3_bit_slice_6534 : p4_bit_slice_6534;
      p5_b <= p5_data_enable ? p4_b : p5_b;
      p5_uge_6502 <= p5_data_enable ? p4_uge_6502 : p5_uge_6502;
      p5_bivisor__1 <= p5_data_enable ? p4_bivisor__1 : p5_bivisor__1;
      p5_uge_6616 <= p5_data_enable ? p4_uge_6616 : p5_uge_6616;
      p5_uge_6694 <= p5_data_enable ? p4_uge_6694 : p5_uge_6694;
      p5_uge_6774 <= p5_data_enable ? p4_uge_6774 : p5_uge_6774;
      p5_uge_6780 <= p5_data_enable ? p4_uge_6780 : p5_uge_6780;
      p5_uge_6858 <= p5_data_enable ? p4_uge_6858 : p5_uge_6858;
      p5_uge_6938 <= p5_data_enable ? uge_6938 : p5_uge_6938;
      p5_r__71 <= p5_data_enable ? r__71 : p5_r__71;
      p5_bit_slice_6510 <= p5_data_enable ? p4_bit_slice_6510 : p5_bit_slice_6510;
      p5_bit_slice_6511 <= p5_data_enable ? p4_bit_slice_6511 : p5_bit_slice_6511;
      p5_bit_slice_6512 <= p5_data_enable ? p4_bit_slice_6512 : p5_bit_slice_6512;
      p5_bit_slice_6513 <= p5_data_enable ? p4_bit_slice_6513 : p5_bit_slice_6513;
      p5_bit_slice_6514 <= p5_data_enable ? p4_bit_slice_6514 : p5_bit_slice_6514;
      p5_bit_slice_6515 <= p5_data_enable ? p4_bit_slice_6515 : p5_bit_slice_6515;
      p5_bit_slice_6516 <= p5_data_enable ? p4_bit_slice_6516 : p5_bit_slice_6516;
      p5_bit_slice_6517 <= p5_data_enable ? p4_bit_slice_6517 : p5_bit_slice_6517;
      p5_bit_slice_6518 <= p5_data_enable ? p4_bit_slice_6518 : p5_bit_slice_6518;
      p5_bit_slice_6519 <= p5_data_enable ? p4_bit_slice_6519 : p5_bit_slice_6519;
      p5_bit_slice_6520 <= p5_data_enable ? p4_bit_slice_6520 : p5_bit_slice_6520;
      p5_bit_slice_6521 <= p5_data_enable ? p4_bit_slice_6521 : p5_bit_slice_6521;
      p5_bit_slice_6522 <= p5_data_enable ? p4_bit_slice_6522 : p5_bit_slice_6522;
      p5_bit_slice_6523 <= p5_data_enable ? p4_bit_slice_6523 : p5_bit_slice_6523;
      p5_bit_slice_6524 <= p5_data_enable ? p4_bit_slice_6524 : p5_bit_slice_6524;
      p5_bit_slice_6525 <= p5_data_enable ? p4_bit_slice_6525 : p5_bit_slice_6525;
      p5_bit_slice_6526 <= p5_data_enable ? p4_bit_slice_6526 : p5_bit_slice_6526;
      p5_bit_slice_6527 <= p5_data_enable ? p4_bit_slice_6527 : p5_bit_slice_6527;
      p5_bit_slice_6528 <= p5_data_enable ? p4_bit_slice_6528 : p5_bit_slice_6528;
      p5_bit_slice_6529 <= p5_data_enable ? p4_bit_slice_6529 : p5_bit_slice_6529;
      p5_bit_slice_6530 <= p5_data_enable ? p4_bit_slice_6530 : p5_bit_slice_6530;
      p5_bit_slice_6531 <= p5_data_enable ? p4_bit_slice_6531 : p5_bit_slice_6531;
      p5_bit_slice_6532 <= p5_data_enable ? p4_bit_slice_6532 : p5_bit_slice_6532;
      p5_bit_slice_6533 <= p5_data_enable ? p4_bit_slice_6533 : p5_bit_slice_6533;
      p5_bit_slice_6534 <= p5_data_enable ? p4_bit_slice_6534 : p5_bit_slice_6534;
      p6_b <= p6_data_enable ? p5_b : p6_b;
      p6_uge_6502 <= p6_data_enable ? p5_uge_6502 : p6_uge_6502;
      p6_bivisor__1 <= p6_data_enable ? p5_bivisor__1 : p6_bivisor__1;
      p6_uge_6616 <= p6_data_enable ? p5_uge_6616 : p6_uge_6616;
      p6_uge_6694 <= p6_data_enable ? p5_uge_6694 : p6_uge_6694;
      p6_uge_6774 <= p6_data_enable ? p5_uge_6774 : p6_uge_6774;
      p6_uge_6780 <= p6_data_enable ? p5_uge_6780 : p6_uge_6780;
      p6_uge_6858 <= p6_data_enable ? p5_uge_6858 : p6_uge_6858;
      p6_uge_6938 <= p6_data_enable ? p5_uge_6938 : p6_uge_6938;
      p6_uge_7016 <= p6_data_enable ? uge_7016 : p6_uge_7016;
      p6_r__72 <= p6_data_enable ? r__72 : p6_r__72;
      p6_bit_slice_6511 <= p6_data_enable ? p5_bit_slice_6511 : p6_bit_slice_6511;
      p6_bit_slice_7019 <= p6_data_enable ? bit_slice_7019 : p6_bit_slice_7019;
      p6_bit_slice_6512 <= p6_data_enable ? p5_bit_slice_6512 : p6_bit_slice_6512;
      p6_bit_slice_6513 <= p6_data_enable ? p5_bit_slice_6513 : p6_bit_slice_6513;
      p6_bit_slice_6514 <= p6_data_enable ? p5_bit_slice_6514 : p6_bit_slice_6514;
      p6_bit_slice_6515 <= p6_data_enable ? p5_bit_slice_6515 : p6_bit_slice_6515;
      p6_bit_slice_6516 <= p6_data_enable ? p5_bit_slice_6516 : p6_bit_slice_6516;
      p6_bit_slice_6517 <= p6_data_enable ? p5_bit_slice_6517 : p6_bit_slice_6517;
      p6_bit_slice_6518 <= p6_data_enable ? p5_bit_slice_6518 : p6_bit_slice_6518;
      p6_bit_slice_6519 <= p6_data_enable ? p5_bit_slice_6519 : p6_bit_slice_6519;
      p6_bit_slice_6520 <= p6_data_enable ? p5_bit_slice_6520 : p6_bit_slice_6520;
      p6_bit_slice_6521 <= p6_data_enable ? p5_bit_slice_6521 : p6_bit_slice_6521;
      p6_bit_slice_6522 <= p6_data_enable ? p5_bit_slice_6522 : p6_bit_slice_6522;
      p6_bit_slice_6523 <= p6_data_enable ? p5_bit_slice_6523 : p6_bit_slice_6523;
      p6_bit_slice_6524 <= p6_data_enable ? p5_bit_slice_6524 : p6_bit_slice_6524;
      p6_bit_slice_6525 <= p6_data_enable ? p5_bit_slice_6525 : p6_bit_slice_6525;
      p6_bit_slice_6526 <= p6_data_enable ? p5_bit_slice_6526 : p6_bit_slice_6526;
      p6_bit_slice_6527 <= p6_data_enable ? p5_bit_slice_6527 : p6_bit_slice_6527;
      p6_bit_slice_6528 <= p6_data_enable ? p5_bit_slice_6528 : p6_bit_slice_6528;
      p6_bit_slice_6529 <= p6_data_enable ? p5_bit_slice_6529 : p6_bit_slice_6529;
      p6_bit_slice_6530 <= p6_data_enable ? p5_bit_slice_6530 : p6_bit_slice_6530;
      p6_bit_slice_6531 <= p6_data_enable ? p5_bit_slice_6531 : p6_bit_slice_6531;
      p6_bit_slice_6532 <= p6_data_enable ? p5_bit_slice_6532 : p6_bit_slice_6532;
      p6_bit_slice_6533 <= p6_data_enable ? p5_bit_slice_6533 : p6_bit_slice_6533;
      p6_bit_slice_6534 <= p6_data_enable ? p5_bit_slice_6534 : p6_bit_slice_6534;
      p7_b <= p7_data_enable ? p6_b : p7_b;
      p7_uge_6502 <= p7_data_enable ? p6_uge_6502 : p7_uge_6502;
      p7_bivisor__1 <= p7_data_enable ? p6_bivisor__1 : p7_bivisor__1;
      p7_uge_6616 <= p7_data_enable ? p6_uge_6616 : p7_uge_6616;
      p7_uge_6694 <= p7_data_enable ? p6_uge_6694 : p7_uge_6694;
      p7_uge_6774 <= p7_data_enable ? p6_uge_6774 : p7_uge_6774;
      p7_uge_6780 <= p7_data_enable ? p6_uge_6780 : p7_uge_6780;
      p7_uge_6858 <= p7_data_enable ? p6_uge_6858 : p7_uge_6858;
      p7_uge_6938 <= p7_data_enable ? p6_uge_6938 : p7_uge_6938;
      p7_uge_7016 <= p7_data_enable ? p6_uge_7016 : p7_uge_7016;
      p7_uge_7096 <= p7_data_enable ? uge_7096 : p7_uge_7096;
      p7_concat_7101 <= p7_data_enable ? concat_7101 : p7_concat_7101;
      p7_uge_7102 <= p7_data_enable ? uge_7102 : p7_uge_7102;
      p7_bit_slice_6513 <= p7_data_enable ? p6_bit_slice_6513 : p7_bit_slice_6513;
      p7_bit_slice_6514 <= p7_data_enable ? p6_bit_slice_6514 : p7_bit_slice_6514;
      p7_bit_slice_6515 <= p7_data_enable ? p6_bit_slice_6515 : p7_bit_slice_6515;
      p7_bit_slice_6516 <= p7_data_enable ? p6_bit_slice_6516 : p7_bit_slice_6516;
      p7_bit_slice_6517 <= p7_data_enable ? p6_bit_slice_6517 : p7_bit_slice_6517;
      p7_bit_slice_6518 <= p7_data_enable ? p6_bit_slice_6518 : p7_bit_slice_6518;
      p7_bit_slice_6519 <= p7_data_enable ? p6_bit_slice_6519 : p7_bit_slice_6519;
      p7_bit_slice_6520 <= p7_data_enable ? p6_bit_slice_6520 : p7_bit_slice_6520;
      p7_bit_slice_6521 <= p7_data_enable ? p6_bit_slice_6521 : p7_bit_slice_6521;
      p7_bit_slice_6522 <= p7_data_enable ? p6_bit_slice_6522 : p7_bit_slice_6522;
      p7_bit_slice_6523 <= p7_data_enable ? p6_bit_slice_6523 : p7_bit_slice_6523;
      p7_bit_slice_6524 <= p7_data_enable ? p6_bit_slice_6524 : p7_bit_slice_6524;
      p7_bit_slice_6525 <= p7_data_enable ? p6_bit_slice_6525 : p7_bit_slice_6525;
      p7_bit_slice_6526 <= p7_data_enable ? p6_bit_slice_6526 : p7_bit_slice_6526;
      p7_bit_slice_6527 <= p7_data_enable ? p6_bit_slice_6527 : p7_bit_slice_6527;
      p7_bit_slice_6528 <= p7_data_enable ? p6_bit_slice_6528 : p7_bit_slice_6528;
      p7_bit_slice_6529 <= p7_data_enable ? p6_bit_slice_6529 : p7_bit_slice_6529;
      p7_bit_slice_6530 <= p7_data_enable ? p6_bit_slice_6530 : p7_bit_slice_6530;
      p7_bit_slice_6531 <= p7_data_enable ? p6_bit_slice_6531 : p7_bit_slice_6531;
      p7_bit_slice_6532 <= p7_data_enable ? p6_bit_slice_6532 : p7_bit_slice_6532;
      p7_bit_slice_6533 <= p7_data_enable ? p6_bit_slice_6533 : p7_bit_slice_6533;
      p7_bit_slice_6534 <= p7_data_enable ? p6_bit_slice_6534 : p7_bit_slice_6534;
      p8_b <= p8_data_enable ? p7_b : p8_b;
      p8_uge_6502 <= p8_data_enable ? p7_uge_6502 : p8_uge_6502;
      p8_bivisor__1 <= p8_data_enable ? p7_bivisor__1 : p8_bivisor__1;
      p8_uge_6616 <= p8_data_enable ? p7_uge_6616 : p8_uge_6616;
      p8_uge_6694 <= p8_data_enable ? p7_uge_6694 : p8_uge_6694;
      p8_uge_6774 <= p8_data_enable ? p7_uge_6774 : p8_uge_6774;
      p8_uge_6780 <= p8_data_enable ? p7_uge_6780 : p8_uge_6780;
      p8_uge_6858 <= p8_data_enable ? p7_uge_6858 : p8_uge_6858;
      p8_uge_6938 <= p8_data_enable ? p7_uge_6938 : p8_uge_6938;
      p8_uge_7016 <= p8_data_enable ? p7_uge_7016 : p8_uge_7016;
      p8_uge_7096 <= p8_data_enable ? p7_uge_7096 : p8_uge_7096;
      p8_uge_7102 <= p8_data_enable ? p7_uge_7102 : p8_uge_7102;
      p8_concat_7179 <= p8_data_enable ? concat_7179 : p8_concat_7179;
      p8_uge_7180 <= p8_data_enable ? uge_7180 : p8_uge_7180;
      p8_sub_7181 <= p8_data_enable ? sub_7181 : p8_sub_7181;
      p8_bit_slice_6514 <= p8_data_enable ? p7_bit_slice_6514 : p8_bit_slice_6514;
      p8_bit_slice_6515 <= p8_data_enable ? p7_bit_slice_6515 : p8_bit_slice_6515;
      p8_bit_slice_6516 <= p8_data_enable ? p7_bit_slice_6516 : p8_bit_slice_6516;
      p8_bit_slice_6517 <= p8_data_enable ? p7_bit_slice_6517 : p8_bit_slice_6517;
      p8_bit_slice_6518 <= p8_data_enable ? p7_bit_slice_6518 : p8_bit_slice_6518;
      p8_bit_slice_6519 <= p8_data_enable ? p7_bit_slice_6519 : p8_bit_slice_6519;
      p8_bit_slice_6520 <= p8_data_enable ? p7_bit_slice_6520 : p8_bit_slice_6520;
      p8_bit_slice_6521 <= p8_data_enable ? p7_bit_slice_6521 : p8_bit_slice_6521;
      p8_bit_slice_6522 <= p8_data_enable ? p7_bit_slice_6522 : p8_bit_slice_6522;
      p8_bit_slice_6523 <= p8_data_enable ? p7_bit_slice_6523 : p8_bit_slice_6523;
      p8_bit_slice_6524 <= p8_data_enable ? p7_bit_slice_6524 : p8_bit_slice_6524;
      p8_bit_slice_6525 <= p8_data_enable ? p7_bit_slice_6525 : p8_bit_slice_6525;
      p8_bit_slice_6526 <= p8_data_enable ? p7_bit_slice_6526 : p8_bit_slice_6526;
      p8_bit_slice_6527 <= p8_data_enable ? p7_bit_slice_6527 : p8_bit_slice_6527;
      p8_bit_slice_6528 <= p8_data_enable ? p7_bit_slice_6528 : p8_bit_slice_6528;
      p8_bit_slice_6529 <= p8_data_enable ? p7_bit_slice_6529 : p8_bit_slice_6529;
      p8_bit_slice_6530 <= p8_data_enable ? p7_bit_slice_6530 : p8_bit_slice_6530;
      p8_bit_slice_6531 <= p8_data_enable ? p7_bit_slice_6531 : p8_bit_slice_6531;
      p8_bit_slice_6532 <= p8_data_enable ? p7_bit_slice_6532 : p8_bit_slice_6532;
      p8_bit_slice_6533 <= p8_data_enable ? p7_bit_slice_6533 : p8_bit_slice_6533;
      p8_bit_slice_6534 <= p8_data_enable ? p7_bit_slice_6534 : p8_bit_slice_6534;
      p9_b <= p9_data_enable ? p8_b : p9_b;
      p9_uge_6502 <= p9_data_enable ? p8_uge_6502 : p9_uge_6502;
      p9_bivisor__1 <= p9_data_enable ? p8_bivisor__1 : p9_bivisor__1;
      p9_uge_6616 <= p9_data_enable ? p8_uge_6616 : p9_uge_6616;
      p9_uge_6694 <= p9_data_enable ? p8_uge_6694 : p9_uge_6694;
      p9_uge_6774 <= p9_data_enable ? p8_uge_6774 : p9_uge_6774;
      p9_uge_6780 <= p9_data_enable ? p8_uge_6780 : p9_uge_6780;
      p9_uge_6858 <= p9_data_enable ? p8_uge_6858 : p9_uge_6858;
      p9_uge_6938 <= p9_data_enable ? p8_uge_6938 : p9_uge_6938;
      p9_uge_7016 <= p9_data_enable ? p8_uge_7016 : p9_uge_7016;
      p9_uge_7096 <= p9_data_enable ? p8_uge_7096 : p9_uge_7096;
      p9_uge_7102 <= p9_data_enable ? p8_uge_7102 : p9_uge_7102;
      p9_uge_7180 <= p9_data_enable ? p8_uge_7180 : p9_uge_7180;
      p9_uge_7260 <= p9_data_enable ? uge_7260 : p9_uge_7260;
      p9_r__76 <= p9_data_enable ? r__76 : p9_r__76;
      p9_bit_slice_6515 <= p9_data_enable ? p8_bit_slice_6515 : p9_bit_slice_6515;
      p9_bit_slice_6516 <= p9_data_enable ? p8_bit_slice_6516 : p9_bit_slice_6516;
      p9_bit_slice_6517 <= p9_data_enable ? p8_bit_slice_6517 : p9_bit_slice_6517;
      p9_bit_slice_6518 <= p9_data_enable ? p8_bit_slice_6518 : p9_bit_slice_6518;
      p9_bit_slice_6519 <= p9_data_enable ? p8_bit_slice_6519 : p9_bit_slice_6519;
      p9_bit_slice_6520 <= p9_data_enable ? p8_bit_slice_6520 : p9_bit_slice_6520;
      p9_bit_slice_6521 <= p9_data_enable ? p8_bit_slice_6521 : p9_bit_slice_6521;
      p9_bit_slice_6522 <= p9_data_enable ? p8_bit_slice_6522 : p9_bit_slice_6522;
      p9_bit_slice_6523 <= p9_data_enable ? p8_bit_slice_6523 : p9_bit_slice_6523;
      p9_bit_slice_6524 <= p9_data_enable ? p8_bit_slice_6524 : p9_bit_slice_6524;
      p9_bit_slice_6525 <= p9_data_enable ? p8_bit_slice_6525 : p9_bit_slice_6525;
      p9_bit_slice_6526 <= p9_data_enable ? p8_bit_slice_6526 : p9_bit_slice_6526;
      p9_bit_slice_6527 <= p9_data_enable ? p8_bit_slice_6527 : p9_bit_slice_6527;
      p9_bit_slice_6528 <= p9_data_enable ? p8_bit_slice_6528 : p9_bit_slice_6528;
      p9_bit_slice_6529 <= p9_data_enable ? p8_bit_slice_6529 : p9_bit_slice_6529;
      p9_bit_slice_6530 <= p9_data_enable ? p8_bit_slice_6530 : p9_bit_slice_6530;
      p9_bit_slice_6531 <= p9_data_enable ? p8_bit_slice_6531 : p9_bit_slice_6531;
      p9_bit_slice_6532 <= p9_data_enable ? p8_bit_slice_6532 : p9_bit_slice_6532;
      p9_bit_slice_6533 <= p9_data_enable ? p8_bit_slice_6533 : p9_bit_slice_6533;
      p9_bit_slice_6534 <= p9_data_enable ? p8_bit_slice_6534 : p9_bit_slice_6534;
      p10_b <= p10_data_enable ? p9_b : p10_b;
      p10_uge_6502 <= p10_data_enable ? p9_uge_6502 : p10_uge_6502;
      p10_bivisor__1 <= p10_data_enable ? p9_bivisor__1 : p10_bivisor__1;
      p10_uge_6616 <= p10_data_enable ? p9_uge_6616 : p10_uge_6616;
      p10_uge_6694 <= p10_data_enable ? p9_uge_6694 : p10_uge_6694;
      p10_uge_6774 <= p10_data_enable ? p9_uge_6774 : p10_uge_6774;
      p10_uge_6780 <= p10_data_enable ? p9_uge_6780 : p10_uge_6780;
      p10_uge_6858 <= p10_data_enable ? p9_uge_6858 : p10_uge_6858;
      p10_uge_6938 <= p10_data_enable ? p9_uge_6938 : p10_uge_6938;
      p10_uge_7016 <= p10_data_enable ? p9_uge_7016 : p10_uge_7016;
      p10_uge_7096 <= p10_data_enable ? p9_uge_7096 : p10_uge_7096;
      p10_uge_7102 <= p10_data_enable ? p9_uge_7102 : p10_uge_7102;
      p10_uge_7180 <= p10_data_enable ? p9_uge_7180 : p10_uge_7180;
      p10_uge_7260 <= p10_data_enable ? p9_uge_7260 : p10_uge_7260;
      p10_uge_7338 <= p10_data_enable ? uge_7338 : p10_uge_7338;
      p10_r__77 <= p10_data_enable ? r__77 : p10_r__77;
      p10_bit_slice_6516 <= p10_data_enable ? p9_bit_slice_6516 : p10_bit_slice_6516;
      p10_bit_slice_7341 <= p10_data_enable ? bit_slice_7341 : p10_bit_slice_7341;
      p10_bit_slice_6517 <= p10_data_enable ? p9_bit_slice_6517 : p10_bit_slice_6517;
      p10_bit_slice_6518 <= p10_data_enable ? p9_bit_slice_6518 : p10_bit_slice_6518;
      p10_bit_slice_6519 <= p10_data_enable ? p9_bit_slice_6519 : p10_bit_slice_6519;
      p10_bit_slice_6520 <= p10_data_enable ? p9_bit_slice_6520 : p10_bit_slice_6520;
      p10_bit_slice_6521 <= p10_data_enable ? p9_bit_slice_6521 : p10_bit_slice_6521;
      p10_bit_slice_6522 <= p10_data_enable ? p9_bit_slice_6522 : p10_bit_slice_6522;
      p10_bit_slice_6523 <= p10_data_enable ? p9_bit_slice_6523 : p10_bit_slice_6523;
      p10_bit_slice_6524 <= p10_data_enable ? p9_bit_slice_6524 : p10_bit_slice_6524;
      p10_bit_slice_6525 <= p10_data_enable ? p9_bit_slice_6525 : p10_bit_slice_6525;
      p10_bit_slice_6526 <= p10_data_enable ? p9_bit_slice_6526 : p10_bit_slice_6526;
      p10_bit_slice_6527 <= p10_data_enable ? p9_bit_slice_6527 : p10_bit_slice_6527;
      p10_bit_slice_6528 <= p10_data_enable ? p9_bit_slice_6528 : p10_bit_slice_6528;
      p10_bit_slice_6529 <= p10_data_enable ? p9_bit_slice_6529 : p10_bit_slice_6529;
      p10_bit_slice_6530 <= p10_data_enable ? p9_bit_slice_6530 : p10_bit_slice_6530;
      p10_bit_slice_6531 <= p10_data_enable ? p9_bit_slice_6531 : p10_bit_slice_6531;
      p10_bit_slice_6532 <= p10_data_enable ? p9_bit_slice_6532 : p10_bit_slice_6532;
      p10_bit_slice_6533 <= p10_data_enable ? p9_bit_slice_6533 : p10_bit_slice_6533;
      p10_bit_slice_6534 <= p10_data_enable ? p9_bit_slice_6534 : p10_bit_slice_6534;
      p11_b <= p11_data_enable ? p10_b : p11_b;
      p11_uge_6502 <= p11_data_enable ? p10_uge_6502 : p11_uge_6502;
      p11_bivisor__1 <= p11_data_enable ? p10_bivisor__1 : p11_bivisor__1;
      p11_uge_6616 <= p11_data_enable ? p10_uge_6616 : p11_uge_6616;
      p11_uge_6694 <= p11_data_enable ? p10_uge_6694 : p11_uge_6694;
      p11_uge_6774 <= p11_data_enable ? p10_uge_6774 : p11_uge_6774;
      p11_uge_6780 <= p11_data_enable ? p10_uge_6780 : p11_uge_6780;
      p11_uge_6858 <= p11_data_enable ? p10_uge_6858 : p11_uge_6858;
      p11_uge_6938 <= p11_data_enable ? p10_uge_6938 : p11_uge_6938;
      p11_uge_7016 <= p11_data_enable ? p10_uge_7016 : p11_uge_7016;
      p11_uge_7096 <= p11_data_enable ? p10_uge_7096 : p11_uge_7096;
      p11_uge_7102 <= p11_data_enable ? p10_uge_7102 : p11_uge_7102;
      p11_uge_7180 <= p11_data_enable ? p10_uge_7180 : p11_uge_7180;
      p11_uge_7260 <= p11_data_enable ? p10_uge_7260 : p11_uge_7260;
      p11_uge_7338 <= p11_data_enable ? p10_uge_7338 : p11_uge_7338;
      p11_uge_7418 <= p11_data_enable ? uge_7418 : p11_uge_7418;
      p11_concat_7423 <= p11_data_enable ? concat_7423 : p11_concat_7423;
      p11_uge_7424 <= p11_data_enable ? uge_7424 : p11_uge_7424;
      p11_bit_slice_6518 <= p11_data_enable ? p10_bit_slice_6518 : p11_bit_slice_6518;
      p11_bit_slice_6519 <= p11_data_enable ? p10_bit_slice_6519 : p11_bit_slice_6519;
      p11_bit_slice_6520 <= p11_data_enable ? p10_bit_slice_6520 : p11_bit_slice_6520;
      p11_bit_slice_6521 <= p11_data_enable ? p10_bit_slice_6521 : p11_bit_slice_6521;
      p11_bit_slice_6522 <= p11_data_enable ? p10_bit_slice_6522 : p11_bit_slice_6522;
      p11_bit_slice_6523 <= p11_data_enable ? p10_bit_slice_6523 : p11_bit_slice_6523;
      p11_bit_slice_6524 <= p11_data_enable ? p10_bit_slice_6524 : p11_bit_slice_6524;
      p11_bit_slice_6525 <= p11_data_enable ? p10_bit_slice_6525 : p11_bit_slice_6525;
      p11_bit_slice_6526 <= p11_data_enable ? p10_bit_slice_6526 : p11_bit_slice_6526;
      p11_bit_slice_6527 <= p11_data_enable ? p10_bit_slice_6527 : p11_bit_slice_6527;
      p11_bit_slice_6528 <= p11_data_enable ? p10_bit_slice_6528 : p11_bit_slice_6528;
      p11_bit_slice_6529 <= p11_data_enable ? p10_bit_slice_6529 : p11_bit_slice_6529;
      p11_bit_slice_6530 <= p11_data_enable ? p10_bit_slice_6530 : p11_bit_slice_6530;
      p11_bit_slice_6531 <= p11_data_enable ? p10_bit_slice_6531 : p11_bit_slice_6531;
      p11_bit_slice_6532 <= p11_data_enable ? p10_bit_slice_6532 : p11_bit_slice_6532;
      p11_bit_slice_6533 <= p11_data_enable ? p10_bit_slice_6533 : p11_bit_slice_6533;
      p11_bit_slice_6534 <= p11_data_enable ? p10_bit_slice_6534 : p11_bit_slice_6534;
      p12_b <= p12_data_enable ? p11_b : p12_b;
      p12_uge_6502 <= p12_data_enable ? p11_uge_6502 : p12_uge_6502;
      p12_bivisor__1 <= p12_data_enable ? p11_bivisor__1 : p12_bivisor__1;
      p12_uge_6616 <= p12_data_enable ? p11_uge_6616 : p12_uge_6616;
      p12_uge_6694 <= p12_data_enable ? p11_uge_6694 : p12_uge_6694;
      p12_uge_6774 <= p12_data_enable ? p11_uge_6774 : p12_uge_6774;
      p12_uge_6780 <= p12_data_enable ? p11_uge_6780 : p12_uge_6780;
      p12_uge_6858 <= p12_data_enable ? p11_uge_6858 : p12_uge_6858;
      p12_uge_6938 <= p12_data_enable ? p11_uge_6938 : p12_uge_6938;
      p12_uge_7016 <= p12_data_enable ? p11_uge_7016 : p12_uge_7016;
      p12_uge_7096 <= p12_data_enable ? p11_uge_7096 : p12_uge_7096;
      p12_uge_7102 <= p12_data_enable ? p11_uge_7102 : p12_uge_7102;
      p12_uge_7180 <= p12_data_enable ? p11_uge_7180 : p12_uge_7180;
      p12_uge_7260 <= p12_data_enable ? p11_uge_7260 : p12_uge_7260;
      p12_uge_7338 <= p12_data_enable ? p11_uge_7338 : p12_uge_7338;
      p12_uge_7418 <= p12_data_enable ? p11_uge_7418 : p12_uge_7418;
      p12_uge_7424 <= p12_data_enable ? p11_uge_7424 : p12_uge_7424;
      p12_concat_7501 <= p12_data_enable ? concat_7501 : p12_concat_7501;
      p12_uge_7502 <= p12_data_enable ? uge_7502 : p12_uge_7502;
      p12_sub_7503 <= p12_data_enable ? sub_7503 : p12_sub_7503;
      p12_bit_slice_6519 <= p12_data_enable ? p11_bit_slice_6519 : p12_bit_slice_6519;
      p12_bit_slice_6520 <= p12_data_enable ? p11_bit_slice_6520 : p12_bit_slice_6520;
      p12_bit_slice_6521 <= p12_data_enable ? p11_bit_slice_6521 : p12_bit_slice_6521;
      p12_bit_slice_6522 <= p12_data_enable ? p11_bit_slice_6522 : p12_bit_slice_6522;
      p12_bit_slice_6523 <= p12_data_enable ? p11_bit_slice_6523 : p12_bit_slice_6523;
      p12_bit_slice_6524 <= p12_data_enable ? p11_bit_slice_6524 : p12_bit_slice_6524;
      p12_bit_slice_6525 <= p12_data_enable ? p11_bit_slice_6525 : p12_bit_slice_6525;
      p12_bit_slice_6526 <= p12_data_enable ? p11_bit_slice_6526 : p12_bit_slice_6526;
      p12_bit_slice_6527 <= p12_data_enable ? p11_bit_slice_6527 : p12_bit_slice_6527;
      p12_bit_slice_6528 <= p12_data_enable ? p11_bit_slice_6528 : p12_bit_slice_6528;
      p12_bit_slice_6529 <= p12_data_enable ? p11_bit_slice_6529 : p12_bit_slice_6529;
      p12_bit_slice_6530 <= p12_data_enable ? p11_bit_slice_6530 : p12_bit_slice_6530;
      p12_bit_slice_6531 <= p12_data_enable ? p11_bit_slice_6531 : p12_bit_slice_6531;
      p12_bit_slice_6532 <= p12_data_enable ? p11_bit_slice_6532 : p12_bit_slice_6532;
      p12_bit_slice_6533 <= p12_data_enable ? p11_bit_slice_6533 : p12_bit_slice_6533;
      p12_bit_slice_6534 <= p12_data_enable ? p11_bit_slice_6534 : p12_bit_slice_6534;
      p13_b <= p13_data_enable ? p12_b : p13_b;
      p13_uge_6502 <= p13_data_enable ? p12_uge_6502 : p13_uge_6502;
      p13_bivisor__1 <= p13_data_enable ? p12_bivisor__1 : p13_bivisor__1;
      p13_uge_6616 <= p13_data_enable ? p12_uge_6616 : p13_uge_6616;
      p13_uge_6694 <= p13_data_enable ? p12_uge_6694 : p13_uge_6694;
      p13_uge_6774 <= p13_data_enable ? p12_uge_6774 : p13_uge_6774;
      p13_uge_6780 <= p13_data_enable ? p12_uge_6780 : p13_uge_6780;
      p13_uge_6858 <= p13_data_enable ? p12_uge_6858 : p13_uge_6858;
      p13_uge_6938 <= p13_data_enable ? p12_uge_6938 : p13_uge_6938;
      p13_uge_7016 <= p13_data_enable ? p12_uge_7016 : p13_uge_7016;
      p13_uge_7096 <= p13_data_enable ? p12_uge_7096 : p13_uge_7096;
      p13_uge_7102 <= p13_data_enable ? p12_uge_7102 : p13_uge_7102;
      p13_uge_7180 <= p13_data_enable ? p12_uge_7180 : p13_uge_7180;
      p13_uge_7260 <= p13_data_enable ? p12_uge_7260 : p13_uge_7260;
      p13_uge_7338 <= p13_data_enable ? p12_uge_7338 : p13_uge_7338;
      p13_uge_7418 <= p13_data_enable ? p12_uge_7418 : p13_uge_7418;
      p13_uge_7424 <= p13_data_enable ? p12_uge_7424 : p13_uge_7424;
      p13_uge_7502 <= p13_data_enable ? p12_uge_7502 : p13_uge_7502;
      p13_uge_7582 <= p13_data_enable ? uge_7582 : p13_uge_7582;
      p13_r__81 <= p13_data_enable ? r__81 : p13_r__81;
      p13_bit_slice_6520 <= p13_data_enable ? p12_bit_slice_6520 : p13_bit_slice_6520;
      p13_bit_slice_6521 <= p13_data_enable ? p12_bit_slice_6521 : p13_bit_slice_6521;
      p13_bit_slice_6522 <= p13_data_enable ? p12_bit_slice_6522 : p13_bit_slice_6522;
      p13_bit_slice_6523 <= p13_data_enable ? p12_bit_slice_6523 : p13_bit_slice_6523;
      p13_bit_slice_6524 <= p13_data_enable ? p12_bit_slice_6524 : p13_bit_slice_6524;
      p13_bit_slice_6525 <= p13_data_enable ? p12_bit_slice_6525 : p13_bit_slice_6525;
      p13_bit_slice_6526 <= p13_data_enable ? p12_bit_slice_6526 : p13_bit_slice_6526;
      p13_bit_slice_6527 <= p13_data_enable ? p12_bit_slice_6527 : p13_bit_slice_6527;
      p13_bit_slice_6528 <= p13_data_enable ? p12_bit_slice_6528 : p13_bit_slice_6528;
      p13_bit_slice_6529 <= p13_data_enable ? p12_bit_slice_6529 : p13_bit_slice_6529;
      p13_bit_slice_6530 <= p13_data_enable ? p12_bit_slice_6530 : p13_bit_slice_6530;
      p13_bit_slice_6531 <= p13_data_enable ? p12_bit_slice_6531 : p13_bit_slice_6531;
      p13_bit_slice_6532 <= p13_data_enable ? p12_bit_slice_6532 : p13_bit_slice_6532;
      p13_bit_slice_6533 <= p13_data_enable ? p12_bit_slice_6533 : p13_bit_slice_6533;
      p13_bit_slice_6534 <= p13_data_enable ? p12_bit_slice_6534 : p13_bit_slice_6534;
      p14_b <= p14_data_enable ? p13_b : p14_b;
      p14_uge_6502 <= p14_data_enable ? p13_uge_6502 : p14_uge_6502;
      p14_bivisor__1 <= p14_data_enable ? p13_bivisor__1 : p14_bivisor__1;
      p14_uge_6616 <= p14_data_enable ? p13_uge_6616 : p14_uge_6616;
      p14_uge_6694 <= p14_data_enable ? p13_uge_6694 : p14_uge_6694;
      p14_uge_6774 <= p14_data_enable ? p13_uge_6774 : p14_uge_6774;
      p14_uge_6780 <= p14_data_enable ? p13_uge_6780 : p14_uge_6780;
      p14_uge_6858 <= p14_data_enable ? p13_uge_6858 : p14_uge_6858;
      p14_uge_6938 <= p14_data_enable ? p13_uge_6938 : p14_uge_6938;
      p14_uge_7016 <= p14_data_enable ? p13_uge_7016 : p14_uge_7016;
      p14_uge_7096 <= p14_data_enable ? p13_uge_7096 : p14_uge_7096;
      p14_uge_7102 <= p14_data_enable ? p13_uge_7102 : p14_uge_7102;
      p14_uge_7180 <= p14_data_enable ? p13_uge_7180 : p14_uge_7180;
      p14_uge_7260 <= p14_data_enable ? p13_uge_7260 : p14_uge_7260;
      p14_uge_7338 <= p14_data_enable ? p13_uge_7338 : p14_uge_7338;
      p14_uge_7418 <= p14_data_enable ? p13_uge_7418 : p14_uge_7418;
      p14_uge_7424 <= p14_data_enable ? p13_uge_7424 : p14_uge_7424;
      p14_uge_7502 <= p14_data_enable ? p13_uge_7502 : p14_uge_7502;
      p14_uge_7582 <= p14_data_enable ? p13_uge_7582 : p14_uge_7582;
      p14_uge_7660 <= p14_data_enable ? uge_7660 : p14_uge_7660;
      p14_r__82 <= p14_data_enable ? r__82 : p14_r__82;
      p14_bit_slice_6521 <= p14_data_enable ? p13_bit_slice_6521 : p14_bit_slice_6521;
      p14_bit_slice_7663 <= p14_data_enable ? bit_slice_7663 : p14_bit_slice_7663;
      p14_bit_slice_6522 <= p14_data_enable ? p13_bit_slice_6522 : p14_bit_slice_6522;
      p14_bit_slice_6523 <= p14_data_enable ? p13_bit_slice_6523 : p14_bit_slice_6523;
      p14_bit_slice_6524 <= p14_data_enable ? p13_bit_slice_6524 : p14_bit_slice_6524;
      p14_bit_slice_6525 <= p14_data_enable ? p13_bit_slice_6525 : p14_bit_slice_6525;
      p14_bit_slice_6526 <= p14_data_enable ? p13_bit_slice_6526 : p14_bit_slice_6526;
      p14_bit_slice_6527 <= p14_data_enable ? p13_bit_slice_6527 : p14_bit_slice_6527;
      p14_bit_slice_6528 <= p14_data_enable ? p13_bit_slice_6528 : p14_bit_slice_6528;
      p14_bit_slice_6529 <= p14_data_enable ? p13_bit_slice_6529 : p14_bit_slice_6529;
      p14_bit_slice_6530 <= p14_data_enable ? p13_bit_slice_6530 : p14_bit_slice_6530;
      p14_bit_slice_6531 <= p14_data_enable ? p13_bit_slice_6531 : p14_bit_slice_6531;
      p14_bit_slice_6532 <= p14_data_enable ? p13_bit_slice_6532 : p14_bit_slice_6532;
      p14_bit_slice_6533 <= p14_data_enable ? p13_bit_slice_6533 : p14_bit_slice_6533;
      p14_bit_slice_6534 <= p14_data_enable ? p13_bit_slice_6534 : p14_bit_slice_6534;
      p15_b <= p15_data_enable ? p14_b : p15_b;
      p15_uge_6502 <= p15_data_enable ? p14_uge_6502 : p15_uge_6502;
      p15_bivisor__1 <= p15_data_enable ? p14_bivisor__1 : p15_bivisor__1;
      p15_uge_6616 <= p15_data_enable ? p14_uge_6616 : p15_uge_6616;
      p15_uge_6694 <= p15_data_enable ? p14_uge_6694 : p15_uge_6694;
      p15_uge_6774 <= p15_data_enable ? p14_uge_6774 : p15_uge_6774;
      p15_uge_6780 <= p15_data_enable ? p14_uge_6780 : p15_uge_6780;
      p15_uge_6858 <= p15_data_enable ? p14_uge_6858 : p15_uge_6858;
      p15_uge_6938 <= p15_data_enable ? p14_uge_6938 : p15_uge_6938;
      p15_uge_7016 <= p15_data_enable ? p14_uge_7016 : p15_uge_7016;
      p15_uge_7096 <= p15_data_enable ? p14_uge_7096 : p15_uge_7096;
      p15_uge_7102 <= p15_data_enable ? p14_uge_7102 : p15_uge_7102;
      p15_uge_7180 <= p15_data_enable ? p14_uge_7180 : p15_uge_7180;
      p15_uge_7260 <= p15_data_enable ? p14_uge_7260 : p15_uge_7260;
      p15_uge_7338 <= p15_data_enable ? p14_uge_7338 : p15_uge_7338;
      p15_uge_7418 <= p15_data_enable ? p14_uge_7418 : p15_uge_7418;
      p15_uge_7424 <= p15_data_enable ? p14_uge_7424 : p15_uge_7424;
      p15_uge_7502 <= p15_data_enable ? p14_uge_7502 : p15_uge_7502;
      p15_uge_7582 <= p15_data_enable ? p14_uge_7582 : p15_uge_7582;
      p15_uge_7660 <= p15_data_enable ? p14_uge_7660 : p15_uge_7660;
      p15_uge_7740 <= p15_data_enable ? uge_7740 : p15_uge_7740;
      p15_concat_7745 <= p15_data_enable ? concat_7745 : p15_concat_7745;
      p15_uge_7746 <= p15_data_enable ? uge_7746 : p15_uge_7746;
      p15_bit_slice_6523 <= p15_data_enable ? p14_bit_slice_6523 : p15_bit_slice_6523;
      p15_bit_slice_6524 <= p15_data_enable ? p14_bit_slice_6524 : p15_bit_slice_6524;
      p15_bit_slice_6525 <= p15_data_enable ? p14_bit_slice_6525 : p15_bit_slice_6525;
      p15_bit_slice_6526 <= p15_data_enable ? p14_bit_slice_6526 : p15_bit_slice_6526;
      p15_bit_slice_6527 <= p15_data_enable ? p14_bit_slice_6527 : p15_bit_slice_6527;
      p15_bit_slice_6528 <= p15_data_enable ? p14_bit_slice_6528 : p15_bit_slice_6528;
      p15_bit_slice_6529 <= p15_data_enable ? p14_bit_slice_6529 : p15_bit_slice_6529;
      p15_bit_slice_6530 <= p15_data_enable ? p14_bit_slice_6530 : p15_bit_slice_6530;
      p15_bit_slice_6531 <= p15_data_enable ? p14_bit_slice_6531 : p15_bit_slice_6531;
      p15_bit_slice_6532 <= p15_data_enable ? p14_bit_slice_6532 : p15_bit_slice_6532;
      p15_bit_slice_6533 <= p15_data_enable ? p14_bit_slice_6533 : p15_bit_slice_6533;
      p15_bit_slice_6534 <= p15_data_enable ? p14_bit_slice_6534 : p15_bit_slice_6534;
      p16_b <= p16_data_enable ? p15_b : p16_b;
      p16_uge_6502 <= p16_data_enable ? p15_uge_6502 : p16_uge_6502;
      p16_bivisor__1 <= p16_data_enable ? p15_bivisor__1 : p16_bivisor__1;
      p16_uge_6616 <= p16_data_enable ? p15_uge_6616 : p16_uge_6616;
      p16_uge_6694 <= p16_data_enable ? p15_uge_6694 : p16_uge_6694;
      p16_uge_6774 <= p16_data_enable ? p15_uge_6774 : p16_uge_6774;
      p16_uge_6780 <= p16_data_enable ? p15_uge_6780 : p16_uge_6780;
      p16_uge_6858 <= p16_data_enable ? p15_uge_6858 : p16_uge_6858;
      p16_uge_6938 <= p16_data_enable ? p15_uge_6938 : p16_uge_6938;
      p16_uge_7016 <= p16_data_enable ? p15_uge_7016 : p16_uge_7016;
      p16_uge_7096 <= p16_data_enable ? p15_uge_7096 : p16_uge_7096;
      p16_uge_7102 <= p16_data_enable ? p15_uge_7102 : p16_uge_7102;
      p16_uge_7180 <= p16_data_enable ? p15_uge_7180 : p16_uge_7180;
      p16_uge_7260 <= p16_data_enable ? p15_uge_7260 : p16_uge_7260;
      p16_uge_7338 <= p16_data_enable ? p15_uge_7338 : p16_uge_7338;
      p16_uge_7418 <= p16_data_enable ? p15_uge_7418 : p16_uge_7418;
      p16_uge_7424 <= p16_data_enable ? p15_uge_7424 : p16_uge_7424;
      p16_uge_7502 <= p16_data_enable ? p15_uge_7502 : p16_uge_7502;
      p16_uge_7582 <= p16_data_enable ? p15_uge_7582 : p16_uge_7582;
      p16_uge_7660 <= p16_data_enable ? p15_uge_7660 : p16_uge_7660;
      p16_uge_7740 <= p16_data_enable ? p15_uge_7740 : p16_uge_7740;
      p16_uge_7746 <= p16_data_enable ? p15_uge_7746 : p16_uge_7746;
      p16_concat_7823 <= p16_data_enable ? concat_7823 : p16_concat_7823;
      p16_uge_7824 <= p16_data_enable ? uge_7824 : p16_uge_7824;
      p16_sub_7825 <= p16_data_enable ? sub_7825 : p16_sub_7825;
      p16_bit_slice_6524 <= p16_data_enable ? p15_bit_slice_6524 : p16_bit_slice_6524;
      p16_bit_slice_6525 <= p16_data_enable ? p15_bit_slice_6525 : p16_bit_slice_6525;
      p16_bit_slice_6526 <= p16_data_enable ? p15_bit_slice_6526 : p16_bit_slice_6526;
      p16_bit_slice_6527 <= p16_data_enable ? p15_bit_slice_6527 : p16_bit_slice_6527;
      p16_bit_slice_6528 <= p16_data_enable ? p15_bit_slice_6528 : p16_bit_slice_6528;
      p16_bit_slice_6529 <= p16_data_enable ? p15_bit_slice_6529 : p16_bit_slice_6529;
      p16_bit_slice_6530 <= p16_data_enable ? p15_bit_slice_6530 : p16_bit_slice_6530;
      p16_bit_slice_6531 <= p16_data_enable ? p15_bit_slice_6531 : p16_bit_slice_6531;
      p16_bit_slice_6532 <= p16_data_enable ? p15_bit_slice_6532 : p16_bit_slice_6532;
      p16_bit_slice_6533 <= p16_data_enable ? p15_bit_slice_6533 : p16_bit_slice_6533;
      p16_bit_slice_6534 <= p16_data_enable ? p15_bit_slice_6534 : p16_bit_slice_6534;
      p17_b <= p17_data_enable ? p16_b : p17_b;
      p17_uge_6502 <= p17_data_enable ? p16_uge_6502 : p17_uge_6502;
      p17_bivisor__1 <= p17_data_enable ? p16_bivisor__1 : p17_bivisor__1;
      p17_uge_6616 <= p17_data_enable ? p16_uge_6616 : p17_uge_6616;
      p17_uge_6694 <= p17_data_enable ? p16_uge_6694 : p17_uge_6694;
      p17_uge_6774 <= p17_data_enable ? p16_uge_6774 : p17_uge_6774;
      p17_uge_6780 <= p17_data_enable ? p16_uge_6780 : p17_uge_6780;
      p17_uge_6858 <= p17_data_enable ? p16_uge_6858 : p17_uge_6858;
      p17_uge_6938 <= p17_data_enable ? p16_uge_6938 : p17_uge_6938;
      p17_uge_7016 <= p17_data_enable ? p16_uge_7016 : p17_uge_7016;
      p17_uge_7096 <= p17_data_enable ? p16_uge_7096 : p17_uge_7096;
      p17_uge_7102 <= p17_data_enable ? p16_uge_7102 : p17_uge_7102;
      p17_uge_7180 <= p17_data_enable ? p16_uge_7180 : p17_uge_7180;
      p17_uge_7260 <= p17_data_enable ? p16_uge_7260 : p17_uge_7260;
      p17_uge_7338 <= p17_data_enable ? p16_uge_7338 : p17_uge_7338;
      p17_uge_7418 <= p17_data_enable ? p16_uge_7418 : p17_uge_7418;
      p17_uge_7424 <= p17_data_enable ? p16_uge_7424 : p17_uge_7424;
      p17_uge_7502 <= p17_data_enable ? p16_uge_7502 : p17_uge_7502;
      p17_uge_7582 <= p17_data_enable ? p16_uge_7582 : p17_uge_7582;
      p17_uge_7660 <= p17_data_enable ? p16_uge_7660 : p17_uge_7660;
      p17_uge_7740 <= p17_data_enable ? p16_uge_7740 : p17_uge_7740;
      p17_uge_7746 <= p17_data_enable ? p16_uge_7746 : p17_uge_7746;
      p17_uge_7824 <= p17_data_enable ? p16_uge_7824 : p17_uge_7824;
      p17_uge_7904 <= p17_data_enable ? uge_7904 : p17_uge_7904;
      p17_r__86 <= p17_data_enable ? r__86 : p17_r__86;
      p17_bit_slice_6525 <= p17_data_enable ? p16_bit_slice_6525 : p17_bit_slice_6525;
      p17_bit_slice_6526 <= p17_data_enable ? p16_bit_slice_6526 : p17_bit_slice_6526;
      p17_bit_slice_6527 <= p17_data_enable ? p16_bit_slice_6527 : p17_bit_slice_6527;
      p17_bit_slice_6528 <= p17_data_enable ? p16_bit_slice_6528 : p17_bit_slice_6528;
      p17_bit_slice_6529 <= p17_data_enable ? p16_bit_slice_6529 : p17_bit_slice_6529;
      p17_bit_slice_6530 <= p17_data_enable ? p16_bit_slice_6530 : p17_bit_slice_6530;
      p17_bit_slice_6531 <= p17_data_enable ? p16_bit_slice_6531 : p17_bit_slice_6531;
      p17_bit_slice_6532 <= p17_data_enable ? p16_bit_slice_6532 : p17_bit_slice_6532;
      p17_bit_slice_6533 <= p17_data_enable ? p16_bit_slice_6533 : p17_bit_slice_6533;
      p17_bit_slice_6534 <= p17_data_enable ? p16_bit_slice_6534 : p17_bit_slice_6534;
      p18_b <= p18_data_enable ? p17_b : p18_b;
      p18_uge_6502 <= p18_data_enable ? p17_uge_6502 : p18_uge_6502;
      p18_bivisor__1 <= p18_data_enable ? p17_bivisor__1 : p18_bivisor__1;
      p18_uge_6616 <= p18_data_enable ? p17_uge_6616 : p18_uge_6616;
      p18_uge_6694 <= p18_data_enable ? p17_uge_6694 : p18_uge_6694;
      p18_uge_6774 <= p18_data_enable ? p17_uge_6774 : p18_uge_6774;
      p18_uge_6780 <= p18_data_enable ? p17_uge_6780 : p18_uge_6780;
      p18_uge_6858 <= p18_data_enable ? p17_uge_6858 : p18_uge_6858;
      p18_uge_6938 <= p18_data_enable ? p17_uge_6938 : p18_uge_6938;
      p18_uge_7016 <= p18_data_enable ? p17_uge_7016 : p18_uge_7016;
      p18_uge_7096 <= p18_data_enable ? p17_uge_7096 : p18_uge_7096;
      p18_uge_7102 <= p18_data_enable ? p17_uge_7102 : p18_uge_7102;
      p18_uge_7180 <= p18_data_enable ? p17_uge_7180 : p18_uge_7180;
      p18_uge_7260 <= p18_data_enable ? p17_uge_7260 : p18_uge_7260;
      p18_uge_7338 <= p18_data_enable ? p17_uge_7338 : p18_uge_7338;
      p18_uge_7418 <= p18_data_enable ? p17_uge_7418 : p18_uge_7418;
      p18_uge_7424 <= p18_data_enable ? p17_uge_7424 : p18_uge_7424;
      p18_uge_7502 <= p18_data_enable ? p17_uge_7502 : p18_uge_7502;
      p18_uge_7582 <= p18_data_enable ? p17_uge_7582 : p18_uge_7582;
      p18_uge_7660 <= p18_data_enable ? p17_uge_7660 : p18_uge_7660;
      p18_uge_7740 <= p18_data_enable ? p17_uge_7740 : p18_uge_7740;
      p18_uge_7746 <= p18_data_enable ? p17_uge_7746 : p18_uge_7746;
      p18_uge_7824 <= p18_data_enable ? p17_uge_7824 : p18_uge_7824;
      p18_uge_7904 <= p18_data_enable ? p17_uge_7904 : p18_uge_7904;
      p18_uge_7982 <= p18_data_enable ? uge_7982 : p18_uge_7982;
      p18_r__87 <= p18_data_enable ? r__87 : p18_r__87;
      p18_bit_slice_6526 <= p18_data_enable ? p17_bit_slice_6526 : p18_bit_slice_6526;
      p18_bit_slice_7985 <= p18_data_enable ? bit_slice_7985 : p18_bit_slice_7985;
      p18_bit_slice_6527 <= p18_data_enable ? p17_bit_slice_6527 : p18_bit_slice_6527;
      p18_bit_slice_6528 <= p18_data_enable ? p17_bit_slice_6528 : p18_bit_slice_6528;
      p18_bit_slice_6529 <= p18_data_enable ? p17_bit_slice_6529 : p18_bit_slice_6529;
      p18_bit_slice_6530 <= p18_data_enable ? p17_bit_slice_6530 : p18_bit_slice_6530;
      p18_bit_slice_6531 <= p18_data_enable ? p17_bit_slice_6531 : p18_bit_slice_6531;
      p18_bit_slice_6532 <= p18_data_enable ? p17_bit_slice_6532 : p18_bit_slice_6532;
      p18_bit_slice_6533 <= p18_data_enable ? p17_bit_slice_6533 : p18_bit_slice_6533;
      p18_bit_slice_6534 <= p18_data_enable ? p17_bit_slice_6534 : p18_bit_slice_6534;
      p19_b <= p19_data_enable ? p18_b : p19_b;
      p19_uge_6502 <= p19_data_enable ? p18_uge_6502 : p19_uge_6502;
      p19_bivisor__1 <= p19_data_enable ? p18_bivisor__1 : p19_bivisor__1;
      p19_uge_6616 <= p19_data_enable ? p18_uge_6616 : p19_uge_6616;
      p19_uge_6694 <= p19_data_enable ? p18_uge_6694 : p19_uge_6694;
      p19_uge_6774 <= p19_data_enable ? p18_uge_6774 : p19_uge_6774;
      p19_uge_6780 <= p19_data_enable ? p18_uge_6780 : p19_uge_6780;
      p19_uge_6858 <= p19_data_enable ? p18_uge_6858 : p19_uge_6858;
      p19_uge_6938 <= p19_data_enable ? p18_uge_6938 : p19_uge_6938;
      p19_uge_7016 <= p19_data_enable ? p18_uge_7016 : p19_uge_7016;
      p19_uge_7096 <= p19_data_enable ? p18_uge_7096 : p19_uge_7096;
      p19_uge_7102 <= p19_data_enable ? p18_uge_7102 : p19_uge_7102;
      p19_uge_7180 <= p19_data_enable ? p18_uge_7180 : p19_uge_7180;
      p19_uge_7260 <= p19_data_enable ? p18_uge_7260 : p19_uge_7260;
      p19_uge_7338 <= p19_data_enable ? p18_uge_7338 : p19_uge_7338;
      p19_uge_7418 <= p19_data_enable ? p18_uge_7418 : p19_uge_7418;
      p19_uge_7424 <= p19_data_enable ? p18_uge_7424 : p19_uge_7424;
      p19_uge_7502 <= p19_data_enable ? p18_uge_7502 : p19_uge_7502;
      p19_uge_7582 <= p19_data_enable ? p18_uge_7582 : p19_uge_7582;
      p19_uge_7660 <= p19_data_enable ? p18_uge_7660 : p19_uge_7660;
      p19_uge_7740 <= p19_data_enable ? p18_uge_7740 : p19_uge_7740;
      p19_uge_7746 <= p19_data_enable ? p18_uge_7746 : p19_uge_7746;
      p19_uge_7824 <= p19_data_enable ? p18_uge_7824 : p19_uge_7824;
      p19_uge_7904 <= p19_data_enable ? p18_uge_7904 : p19_uge_7904;
      p19_uge_7982 <= p19_data_enable ? p18_uge_7982 : p19_uge_7982;
      p19_uge_8062 <= p19_data_enable ? uge_8062 : p19_uge_8062;
      p19_concat_8067 <= p19_data_enable ? concat_8067 : p19_concat_8067;
      p19_uge_8068 <= p19_data_enable ? uge_8068 : p19_uge_8068;
      p19_bit_slice_6528 <= p19_data_enable ? p18_bit_slice_6528 : p19_bit_slice_6528;
      p19_bit_slice_6529 <= p19_data_enable ? p18_bit_slice_6529 : p19_bit_slice_6529;
      p19_bit_slice_6530 <= p19_data_enable ? p18_bit_slice_6530 : p19_bit_slice_6530;
      p19_bit_slice_6531 <= p19_data_enable ? p18_bit_slice_6531 : p19_bit_slice_6531;
      p19_bit_slice_6532 <= p19_data_enable ? p18_bit_slice_6532 : p19_bit_slice_6532;
      p19_bit_slice_6533 <= p19_data_enable ? p18_bit_slice_6533 : p19_bit_slice_6533;
      p19_bit_slice_6534 <= p19_data_enable ? p18_bit_slice_6534 : p19_bit_slice_6534;
      p20_b <= p20_data_enable ? p19_b : p20_b;
      p20_uge_6502 <= p20_data_enable ? p19_uge_6502 : p20_uge_6502;
      p20_bivisor__1 <= p20_data_enable ? p19_bivisor__1 : p20_bivisor__1;
      p20_uge_6616 <= p20_data_enable ? p19_uge_6616 : p20_uge_6616;
      p20_uge_6694 <= p20_data_enable ? p19_uge_6694 : p20_uge_6694;
      p20_uge_6774 <= p20_data_enable ? p19_uge_6774 : p20_uge_6774;
      p20_uge_6780 <= p20_data_enable ? p19_uge_6780 : p20_uge_6780;
      p20_uge_6858 <= p20_data_enable ? p19_uge_6858 : p20_uge_6858;
      p20_uge_6938 <= p20_data_enable ? p19_uge_6938 : p20_uge_6938;
      p20_uge_7016 <= p20_data_enable ? p19_uge_7016 : p20_uge_7016;
      p20_uge_7096 <= p20_data_enable ? p19_uge_7096 : p20_uge_7096;
      p20_uge_7102 <= p20_data_enable ? p19_uge_7102 : p20_uge_7102;
      p20_uge_7180 <= p20_data_enable ? p19_uge_7180 : p20_uge_7180;
      p20_uge_7260 <= p20_data_enable ? p19_uge_7260 : p20_uge_7260;
      p20_uge_7338 <= p20_data_enable ? p19_uge_7338 : p20_uge_7338;
      p20_uge_7418 <= p20_data_enable ? p19_uge_7418 : p20_uge_7418;
      p20_uge_7424 <= p20_data_enable ? p19_uge_7424 : p20_uge_7424;
      p20_uge_7502 <= p20_data_enable ? p19_uge_7502 : p20_uge_7502;
      p20_uge_7582 <= p20_data_enable ? p19_uge_7582 : p20_uge_7582;
      p20_uge_7660 <= p20_data_enable ? p19_uge_7660 : p20_uge_7660;
      p20_uge_7740 <= p20_data_enable ? p19_uge_7740 : p20_uge_7740;
      p20_uge_7746 <= p20_data_enable ? p19_uge_7746 : p20_uge_7746;
      p20_uge_7824 <= p20_data_enable ? p19_uge_7824 : p20_uge_7824;
      p20_uge_7904 <= p20_data_enable ? p19_uge_7904 : p20_uge_7904;
      p20_uge_7982 <= p20_data_enable ? p19_uge_7982 : p20_uge_7982;
      p20_uge_8062 <= p20_data_enable ? p19_uge_8062 : p20_uge_8062;
      p20_uge_8068 <= p20_data_enable ? p19_uge_8068 : p20_uge_8068;
      p20_concat_8145 <= p20_data_enable ? concat_8145 : p20_concat_8145;
      p20_uge_8146 <= p20_data_enable ? uge_8146 : p20_uge_8146;
      p20_sub_8147 <= p20_data_enable ? sub_8147 : p20_sub_8147;
      p20_bit_slice_6529 <= p20_data_enable ? p19_bit_slice_6529 : p20_bit_slice_6529;
      p20_bit_slice_6530 <= p20_data_enable ? p19_bit_slice_6530 : p20_bit_slice_6530;
      p20_bit_slice_6531 <= p20_data_enable ? p19_bit_slice_6531 : p20_bit_slice_6531;
      p20_bit_slice_6532 <= p20_data_enable ? p19_bit_slice_6532 : p20_bit_slice_6532;
      p20_bit_slice_6533 <= p20_data_enable ? p19_bit_slice_6533 : p20_bit_slice_6533;
      p20_bit_slice_6534 <= p20_data_enable ? p19_bit_slice_6534 : p20_bit_slice_6534;
      p21_b <= p21_data_enable ? p20_b : p21_b;
      p21_uge_6502 <= p21_data_enable ? p20_uge_6502 : p21_uge_6502;
      p21_bivisor__1 <= p21_data_enable ? p20_bivisor__1 : p21_bivisor__1;
      p21_uge_6616 <= p21_data_enable ? p20_uge_6616 : p21_uge_6616;
      p21_uge_6694 <= p21_data_enable ? p20_uge_6694 : p21_uge_6694;
      p21_uge_6774 <= p21_data_enable ? p20_uge_6774 : p21_uge_6774;
      p21_uge_6780 <= p21_data_enable ? p20_uge_6780 : p21_uge_6780;
      p21_uge_6858 <= p21_data_enable ? p20_uge_6858 : p21_uge_6858;
      p21_uge_6938 <= p21_data_enable ? p20_uge_6938 : p21_uge_6938;
      p21_uge_7016 <= p21_data_enable ? p20_uge_7016 : p21_uge_7016;
      p21_uge_7096 <= p21_data_enable ? p20_uge_7096 : p21_uge_7096;
      p21_uge_7102 <= p21_data_enable ? p20_uge_7102 : p21_uge_7102;
      p21_uge_7180 <= p21_data_enable ? p20_uge_7180 : p21_uge_7180;
      p21_uge_7260 <= p21_data_enable ? p20_uge_7260 : p21_uge_7260;
      p21_uge_7338 <= p21_data_enable ? p20_uge_7338 : p21_uge_7338;
      p21_uge_7418 <= p21_data_enable ? p20_uge_7418 : p21_uge_7418;
      p21_uge_7424 <= p21_data_enable ? p20_uge_7424 : p21_uge_7424;
      p21_uge_7502 <= p21_data_enable ? p20_uge_7502 : p21_uge_7502;
      p21_uge_7582 <= p21_data_enable ? p20_uge_7582 : p21_uge_7582;
      p21_uge_7660 <= p21_data_enable ? p20_uge_7660 : p21_uge_7660;
      p21_uge_7740 <= p21_data_enable ? p20_uge_7740 : p21_uge_7740;
      p21_uge_7746 <= p21_data_enable ? p20_uge_7746 : p21_uge_7746;
      p21_uge_7824 <= p21_data_enable ? p20_uge_7824 : p21_uge_7824;
      p21_uge_7904 <= p21_data_enable ? p20_uge_7904 : p21_uge_7904;
      p21_uge_7982 <= p21_data_enable ? p20_uge_7982 : p21_uge_7982;
      p21_uge_8062 <= p21_data_enable ? p20_uge_8062 : p21_uge_8062;
      p21_uge_8068 <= p21_data_enable ? p20_uge_8068 : p21_uge_8068;
      p21_uge_8146 <= p21_data_enable ? p20_uge_8146 : p21_uge_8146;
      p21_uge_8226 <= p21_data_enable ? uge_8226 : p21_uge_8226;
      p21_r__91 <= p21_data_enable ? r__91 : p21_r__91;
      p21_bit_slice_6530 <= p21_data_enable ? p20_bit_slice_6530 : p21_bit_slice_6530;
      p21_bit_slice_6531 <= p21_data_enable ? p20_bit_slice_6531 : p21_bit_slice_6531;
      p21_bit_slice_6532 <= p21_data_enable ? p20_bit_slice_6532 : p21_bit_slice_6532;
      p21_bit_slice_6533 <= p21_data_enable ? p20_bit_slice_6533 : p21_bit_slice_6533;
      p21_bit_slice_6534 <= p21_data_enable ? p20_bit_slice_6534 : p21_bit_slice_6534;
      p22_b <= p22_data_enable ? p21_b : p22_b;
      p22_uge_6502 <= p22_data_enable ? p21_uge_6502 : p22_uge_6502;
      p22_bivisor__1 <= p22_data_enable ? p21_bivisor__1 : p22_bivisor__1;
      p22_uge_6616 <= p22_data_enable ? p21_uge_6616 : p22_uge_6616;
      p22_uge_6694 <= p22_data_enable ? p21_uge_6694 : p22_uge_6694;
      p22_uge_6774 <= p22_data_enable ? p21_uge_6774 : p22_uge_6774;
      p22_uge_6780 <= p22_data_enable ? p21_uge_6780 : p22_uge_6780;
      p22_uge_6858 <= p22_data_enable ? p21_uge_6858 : p22_uge_6858;
      p22_uge_6938 <= p22_data_enable ? p21_uge_6938 : p22_uge_6938;
      p22_uge_7016 <= p22_data_enable ? p21_uge_7016 : p22_uge_7016;
      p22_uge_7096 <= p22_data_enable ? p21_uge_7096 : p22_uge_7096;
      p22_uge_7102 <= p22_data_enable ? p21_uge_7102 : p22_uge_7102;
      p22_uge_7180 <= p22_data_enable ? p21_uge_7180 : p22_uge_7180;
      p22_uge_7260 <= p22_data_enable ? p21_uge_7260 : p22_uge_7260;
      p22_uge_7338 <= p22_data_enable ? p21_uge_7338 : p22_uge_7338;
      p22_uge_7418 <= p22_data_enable ? p21_uge_7418 : p22_uge_7418;
      p22_uge_7424 <= p22_data_enable ? p21_uge_7424 : p22_uge_7424;
      p22_uge_7502 <= p22_data_enable ? p21_uge_7502 : p22_uge_7502;
      p22_uge_7582 <= p22_data_enable ? p21_uge_7582 : p22_uge_7582;
      p22_uge_7660 <= p22_data_enable ? p21_uge_7660 : p22_uge_7660;
      p22_uge_7740 <= p22_data_enable ? p21_uge_7740 : p22_uge_7740;
      p22_uge_7746 <= p22_data_enable ? p21_uge_7746 : p22_uge_7746;
      p22_uge_7824 <= p22_data_enable ? p21_uge_7824 : p22_uge_7824;
      p22_uge_7904 <= p22_data_enable ? p21_uge_7904 : p22_uge_7904;
      p22_uge_7982 <= p22_data_enable ? p21_uge_7982 : p22_uge_7982;
      p22_uge_8062 <= p22_data_enable ? p21_uge_8062 : p22_uge_8062;
      p22_uge_8068 <= p22_data_enable ? p21_uge_8068 : p22_uge_8068;
      p22_uge_8146 <= p22_data_enable ? p21_uge_8146 : p22_uge_8146;
      p22_uge_8226 <= p22_data_enable ? p21_uge_8226 : p22_uge_8226;
      p22_uge_8304 <= p22_data_enable ? uge_8304 : p22_uge_8304;
      p22_r__92 <= p22_data_enable ? r__92 : p22_r__92;
      p22_bit_slice_6531 <= p22_data_enable ? p21_bit_slice_6531 : p22_bit_slice_6531;
      p22_bit_slice_8307 <= p22_data_enable ? bit_slice_8307 : p22_bit_slice_8307;
      p22_bit_slice_6532 <= p22_data_enable ? p21_bit_slice_6532 : p22_bit_slice_6532;
      p22_bit_slice_6533 <= p22_data_enable ? p21_bit_slice_6533 : p22_bit_slice_6533;
      p22_bit_slice_6534 <= p22_data_enable ? p21_bit_slice_6534 : p22_bit_slice_6534;
      p23_b <= p23_data_enable ? p22_b : p23_b;
      p23_uge_6502 <= p23_data_enable ? p22_uge_6502 : p23_uge_6502;
      p23_bivisor__1 <= p23_data_enable ? p22_bivisor__1 : p23_bivisor__1;
      p23_uge_6616 <= p23_data_enable ? p22_uge_6616 : p23_uge_6616;
      p23_uge_6694 <= p23_data_enable ? p22_uge_6694 : p23_uge_6694;
      p23_uge_6774 <= p23_data_enable ? p22_uge_6774 : p23_uge_6774;
      p23_uge_6780 <= p23_data_enable ? p22_uge_6780 : p23_uge_6780;
      p23_uge_6858 <= p23_data_enable ? p22_uge_6858 : p23_uge_6858;
      p23_uge_6938 <= p23_data_enable ? p22_uge_6938 : p23_uge_6938;
      p23_uge_7016 <= p23_data_enable ? p22_uge_7016 : p23_uge_7016;
      p23_uge_7096 <= p23_data_enable ? p22_uge_7096 : p23_uge_7096;
      p23_uge_7102 <= p23_data_enable ? p22_uge_7102 : p23_uge_7102;
      p23_uge_7180 <= p23_data_enable ? p22_uge_7180 : p23_uge_7180;
      p23_uge_7260 <= p23_data_enable ? p22_uge_7260 : p23_uge_7260;
      p23_uge_7338 <= p23_data_enable ? p22_uge_7338 : p23_uge_7338;
      p23_uge_7418 <= p23_data_enable ? p22_uge_7418 : p23_uge_7418;
      p23_uge_7424 <= p23_data_enable ? p22_uge_7424 : p23_uge_7424;
      p23_uge_7502 <= p23_data_enable ? p22_uge_7502 : p23_uge_7502;
      p23_uge_7582 <= p23_data_enable ? p22_uge_7582 : p23_uge_7582;
      p23_uge_7660 <= p23_data_enable ? p22_uge_7660 : p23_uge_7660;
      p23_uge_7740 <= p23_data_enable ? p22_uge_7740 : p23_uge_7740;
      p23_uge_7746 <= p23_data_enable ? p22_uge_7746 : p23_uge_7746;
      p23_uge_7824 <= p23_data_enable ? p22_uge_7824 : p23_uge_7824;
      p23_uge_7904 <= p23_data_enable ? p22_uge_7904 : p23_uge_7904;
      p23_uge_7982 <= p23_data_enable ? p22_uge_7982 : p23_uge_7982;
      p23_uge_8062 <= p23_data_enable ? p22_uge_8062 : p23_uge_8062;
      p23_uge_8068 <= p23_data_enable ? p22_uge_8068 : p23_uge_8068;
      p23_uge_8146 <= p23_data_enable ? p22_uge_8146 : p23_uge_8146;
      p23_uge_8226 <= p23_data_enable ? p22_uge_8226 : p23_uge_8226;
      p23_uge_8304 <= p23_data_enable ? p22_uge_8304 : p23_uge_8304;
      p23_uge_8384 <= p23_data_enable ? uge_8384 : p23_uge_8384;
      p23_concat_8389 <= p23_data_enable ? concat_8389 : p23_concat_8389;
      p23_uge_8390 <= p23_data_enable ? uge_8390 : p23_uge_8390;
      p23_bit_slice_6533 <= p23_data_enable ? p22_bit_slice_6533 : p23_bit_slice_6533;
      p23_bit_slice_6534 <= p23_data_enable ? p22_bit_slice_6534 : p23_bit_slice_6534;
      p24_uge_6502 <= p24_data_enable ? p23_uge_6502 : p24_uge_6502;
      p24_bivisor__1 <= p24_data_enable ? p23_bivisor__1 : p24_bivisor__1;
      p24_uge_6616 <= p24_data_enable ? p23_uge_6616 : p24_uge_6616;
      p24_uge_6694 <= p24_data_enable ? p23_uge_6694 : p24_uge_6694;
      p24_uge_6774 <= p24_data_enable ? p23_uge_6774 : p24_uge_6774;
      p24_uge_6780 <= p24_data_enable ? p23_uge_6780 : p24_uge_6780;
      p24_uge_6858 <= p24_data_enable ? p23_uge_6858 : p24_uge_6858;
      p24_uge_6938 <= p24_data_enable ? p23_uge_6938 : p24_uge_6938;
      p24_uge_7016 <= p24_data_enable ? p23_uge_7016 : p24_uge_7016;
      p24_uge_7096 <= p24_data_enable ? p23_uge_7096 : p24_uge_7096;
      p24_uge_7102 <= p24_data_enable ? p23_uge_7102 : p24_uge_7102;
      p24_uge_7180 <= p24_data_enable ? p23_uge_7180 : p24_uge_7180;
      p24_uge_7260 <= p24_data_enable ? p23_uge_7260 : p24_uge_7260;
      p24_uge_7338 <= p24_data_enable ? p23_uge_7338 : p24_uge_7338;
      p24_uge_7418 <= p24_data_enable ? p23_uge_7418 : p24_uge_7418;
      p24_uge_7424 <= p24_data_enable ? p23_uge_7424 : p24_uge_7424;
      p24_uge_7502 <= p24_data_enable ? p23_uge_7502 : p24_uge_7502;
      p24_uge_7582 <= p24_data_enable ? p23_uge_7582 : p24_uge_7582;
      p24_uge_7660 <= p24_data_enable ? p23_uge_7660 : p24_uge_7660;
      p24_uge_7740 <= p24_data_enable ? p23_uge_7740 : p24_uge_7740;
      p24_uge_7746 <= p24_data_enable ? p23_uge_7746 : p24_uge_7746;
      p24_uge_7824 <= p24_data_enable ? p23_uge_7824 : p24_uge_7824;
      p24_uge_7904 <= p24_data_enable ? p23_uge_7904 : p24_uge_7904;
      p24_uge_7982 <= p24_data_enable ? p23_uge_7982 : p24_uge_7982;
      p24_uge_8062 <= p24_data_enable ? p23_uge_8062 : p24_uge_8062;
      p24_uge_8068 <= p24_data_enable ? p23_uge_8068 : p24_uge_8068;
      p24_uge_8146 <= p24_data_enable ? p23_uge_8146 : p24_uge_8146;
      p24_uge_8226 <= p24_data_enable ? p23_uge_8226 : p24_uge_8226;
      p24_uge_8304 <= p24_data_enable ? p23_uge_8304 : p24_uge_8304;
      p24_uge_8384 <= p24_data_enable ? p23_uge_8384 : p24_uge_8384;
      p24_uge_8390 <= p24_data_enable ? p23_uge_8390 : p24_uge_8390;
      p24_concat_8467 <= p24_data_enable ? concat_8467 : p24_concat_8467;
      p24_uge_8468 <= p24_data_enable ? uge_8468 : p24_uge_8468;
      p24_sub_8469 <= p24_data_enable ? sub_8469 : p24_sub_8469;
      p24_bit_slice_6534 <= p24_data_enable ? p23_bit_slice_6534 : p24_bit_slice_6534;
      p0_valid <= p0_enable ? p0_all_active_inputs_valid : p0_valid;
      p1_valid <= p1_enable ? p0_valid : p1_valid;
      p2_valid <= p2_enable ? p1_valid : p2_valid;
      p3_valid <= p3_enable ? p2_valid : p3_valid;
      p4_valid <= p4_enable ? p3_valid : p4_valid;
      p5_valid <= p5_enable ? p4_valid : p5_valid;
      p6_valid <= p6_enable ? p5_valid : p6_valid;
      p7_valid <= p7_enable ? p6_valid : p7_valid;
      p8_valid <= p8_enable ? p7_valid : p8_valid;
      p9_valid <= p9_enable ? p8_valid : p9_valid;
      p10_valid <= p10_enable ? p9_valid : p10_valid;
      p11_valid <= p11_enable ? p10_valid : p11_valid;
      p12_valid <= p12_enable ? p11_valid : p12_valid;
      p13_valid <= p13_enable ? p12_valid : p13_valid;
      p14_valid <= p14_enable ? p13_valid : p14_valid;
      p15_valid <= p15_enable ? p14_valid : p15_valid;
      p16_valid <= p16_enable ? p15_valid : p16_valid;
      p17_valid <= p17_enable ? p16_valid : p17_valid;
      p18_valid <= p18_enable ? p17_valid : p18_valid;
      p19_valid <= p19_enable ? p18_valid : p19_valid;
      p20_valid <= p20_enable ? p19_valid : p20_valid;
      p21_valid <= p21_enable ? p20_valid : p21_valid;
      p22_valid <= p22_enable ? p21_valid : p22_valid;
      p23_valid <= p23_enable ? p22_valid : p23_valid;
      p24_valid <= p24_enable ? p23_valid : p24_valid;
      p25_valid <= p25_enable ? p25_stage_done : p25_valid;
      p26_valid <= p26_enable ? p25_valid : p26_valid;
      p27_valid <= p27_enable ? p26_valid : p27_valid;
      p28_valid <= p28_enable ? p27_valid : p28_valid;
      p29_valid <= p29_enable ? p28_valid : p29_valid;
      p30_valid <= p30_enable ? p29_valid : p30_valid;
      lhs_reg <= lhs_load_en ? lhs : lhs_reg;
      lhs_valid_reg <= lhs_valid_load_en ? lhs_valid : lhs_valid_reg;
      rhs_reg <= rhs_load_en ? rhs : rhs_reg;
      rhs_valid_reg <= rhs_valid_load_en ? rhs_valid : rhs_valid_reg;
      result_reg <= result_load_en ? q__32 : result_reg;
      result_valid_reg <= result_valid_load_en ? p24_valid : result_valid_reg;
    end
  end
  assign result = result_reg;
  assign result_valid = result_valid_reg;
  assign lhs_ready = lhs_load_en;
  assign rhs_ready = rhs_load_en;
endmodule
module xls_subf32(
  input wire clk,
  input wire rst,
  input wire [31:0] rhs,
  input wire rhs_valid,
  input wire [31:0] lhs,
  input wire lhs_valid,
  input wire result_ready,
  output wire [31:0] result,
  output wire result_valid,
  output wire rhs_ready,
  output wire lhs_ready
);
  function automatic [3:0] priority_sel_4b_2way (input reg [1:0] sel, input reg [3:0] case0, input reg [3:0] case1, input reg [3:0] default_value);
    begin
      casez (sel)
        2'b?1: begin
          priority_sel_4b_2way = case0;
        end
        2'b10: begin
          priority_sel_4b_2way = case1;
        end
        2'b00: begin
          priority_sel_4b_2way = default_value;
        end
        default: begin
          // Propagate X
          priority_sel_4b_2way = 4'dx;
        end
      endcase
    end
  endfunction
  function automatic [1:0] priority_sel_2b_2way (input reg [1:0] sel, input reg [1:0] case0, input reg [1:0] case1, input reg [1:0] default_value);
    begin
      casez (sel)
        2'b?1: begin
          priority_sel_2b_2way = case0;
        end
        2'b10: begin
          priority_sel_2b_2way = case1;
        end
        2'b00: begin
          priority_sel_2b_2way = default_value;
        end
        default: begin
          // Propagate X
          priority_sel_2b_2way = 2'dx;
        end
      endcase
    end
  endfunction
  function automatic priority_sel_1b_4way (input reg [3:0] sel, input reg case0, input reg case1, input reg case2, input reg case3, input reg default_value);
    begin
      casez (sel)
        4'b???1: begin
          priority_sel_1b_4way = case0;
        end
        4'b??10: begin
          priority_sel_1b_4way = case1;
        end
        4'b?100: begin
          priority_sel_1b_4way = case2;
        end
        4'b1000: begin
          priority_sel_1b_4way = case3;
        end
        4'b0000: begin
          priority_sel_1b_4way = default_value;
        end
        default: begin
          // Propagate X
          priority_sel_1b_4way = 1'dx;
        end
      endcase
    end
  endfunction
  function automatic priority_sel_1b_3way (input reg [2:0] sel, input reg case0, input reg case1, input reg case2, input reg default_value);
    begin
      casez (sel)
        3'b??1: begin
          priority_sel_1b_3way = case0;
        end
        3'b?10: begin
          priority_sel_1b_3way = case1;
        end
        3'b100: begin
          priority_sel_1b_3way = case2;
        end
        3'b000: begin
          priority_sel_1b_3way = default_value;
        end
        default: begin
          // Propagate X
          priority_sel_1b_3way = 1'dx;
        end
      endcase
    end
  endfunction
  function automatic [2:0] priority_sel_3b_2way (input reg [1:0] sel, input reg [2:0] case0, input reg [2:0] case1, input reg [2:0] default_value);
    begin
      casez (sel)
        2'b?1: begin
          priority_sel_3b_2way = case0;
        end
        2'b10: begin
          priority_sel_3b_2way = case1;
        end
        2'b00: begin
          priority_sel_3b_2way = default_value;
        end
        default: begin
          // Propagate X
          priority_sel_3b_2way = 3'dx;
        end
      endcase
    end
  endfunction
  function automatic [1:0] priority_sel_2b_4way (input reg [3:0] sel, input reg [1:0] case0, input reg [1:0] case1, input reg [1:0] case2, input reg [1:0] case3, input reg [1:0] default_value);
    begin
      casez (sel)
        4'b???1: begin
          priority_sel_2b_4way = case0;
        end
        4'b??10: begin
          priority_sel_2b_4way = case1;
        end
        4'b?100: begin
          priority_sel_2b_4way = case2;
        end
        4'b1000: begin
          priority_sel_2b_4way = case3;
        end
        4'b0000: begin
          priority_sel_2b_4way = default_value;
        end
        default: begin
          // Propagate X
          priority_sel_2b_4way = 2'dx;
        end
      endcase
    end
  endfunction
  function automatic priority_sel_1b_2way (input reg [1:0] sel, input reg case0, input reg case1, input reg default_value);
    begin
      casez (sel)
        2'b?1: begin
          priority_sel_1b_2way = case0;
        end
        2'b10: begin
          priority_sel_1b_2way = case1;
        end
        2'b00: begin
          priority_sel_1b_2way = default_value;
        end
        default: begin
          // Propagate X
          priority_sel_1b_2way = 1'dx;
        end
      endcase
    end
  endfunction
  wire [31:0] rhs_reg_init = {1'h0, 8'h00, 23'h00_0000};
  wire [31:0] lhs_reg_init = {1'h0, 8'h00, 23'h00_0000};
  wire [31:0] result_reg_init = {1'h0, 8'h00, 23'h00_0000};
  reg [7:0] p0_b_bexp__4;
  reg [7:0] p0_a_bexp__2;
  reg p0_bit_slice_21156;
  reg [22:0] p0_b_fraction__4;
  reg [22:0] p0_tuple_index_21158;
  reg [7:0] p0_bit_slice_21159;
  reg p0_not_21161;
  reg p0_tuple_index_21162;
  reg [7:0] p1_a_bexp__4;
  reg p1_b_sign__3;
  reg p1_xor_21216;
  reg [24:0] p1_wide_x_squeezed;
  reg [24:0] p1_bit_slice_21218;
  reg [27:0] p1_shrl_21219;
  reg p1_sticky;
  reg p1_is_operand_inf;
  reg p1_and_21249;
  reg p1_is_result_nan;
  reg p1_not_21251;
  reg [7:0] p2_a_bexp__4;
  reg [27:0] p2_abs_fraction__1;
  reg p2_not_21297;
  reg p2_is_operand_inf;
  reg p2_is_result_nan;
  reg p2_result_sign;
  reg p2_not_21251;
  reg [7:0] p3_a_bexp__4;
  reg [27:0] p3_abs_fraction__1;
  reg p3_carry_bit;
  reg p3_and_21438;
  reg p3_and_21440;
  reg p3_nor_21446;
  reg p3_nor_21473;
  reg p3_and_21474;
  reg [2:0] p3_priority_sel_21475;
  reg [1:0] p3_priority_sel_21476;
  reg [2:0] p3_priority_sel_21477;
  reg p3_or_21478;
  reg p3_not_21297;
  reg p3_is_operand_inf;
  reg p3_is_result_nan;
  reg p3_result_sign__2;
  reg [7:0] p4_a_bexp__4;
  reg p4_and_21474;
  reg [3:0] p4_leading_zeroes__0_to_4;
  reg [2:0] p4_normal_chunk;
  reg [1:0] p4_half_way_chunk;
  reg [23:0] p4_bit_slice_21532;
  reg p4_not_21297;
  reg p4_is_operand_inf;
  reg p4_is_result_nan;
  reg p4_result_sign__2;
  reg p5_and_21474;
  reg [3:0] p5_leading_zeroes__0_to_4;
  reg [9:0] p5_concat_21572;
  reg p5_not_21297;
  reg p5_is_operand_inf;
  reg p5_is_result_nan;
  reg [22:0] p5_result_fraction;
  reg p5_result_sign__2;
  reg [8:0] p6_wide_exponent__2;
  reg p6_is_operand_inf;
  reg p6_is_result_nan;
  reg [22:0] p6_result_fraction;
  reg p6_result_sign__2;
  reg p7_is_result_nan;
  reg [22:0] p7_result_fraction__3;
  reg p7_result_sign__2;
  reg [7:0] p7_result_exponent__2;
  reg p0_valid;
  reg p1_valid;
  reg p2_valid;
  reg p3_valid;
  reg p4_valid;
  reg p5_valid;
  reg p6_valid;
  reg p7_valid;
  reg [31:0] rhs_reg;
  reg rhs_valid_reg;
  reg [31:0] lhs_reg;
  reg lhs_valid_reg;
  reg [31:0] result_reg;
  reg result_valid_reg;
  wire result_valid_inv;
  wire result_valid_load_en;
  wire result_load_en;
  wire p8_stage_done;
  wire p8_not_valid;
  wire p7_enable;
  wire p7_data_enable;
  wire p7_not_valid;
  wire p6_enable;
  wire p6_data_enable;
  wire p6_not_valid;
  wire p5_enable;
  wire p5_data_enable;
  wire p5_not_valid;
  wire p4_enable;
  wire p4_data_enable;
  wire p4_not_valid;
  wire p3_enable;
  wire p3_data_enable;
  wire p3_not_valid;
  wire [2:0] fraction_shift__3;
  wire p2_enable;
  wire [9:0] add_21599;
  wire [24:0] concat_21560;
  wire carry_bit;
  wire [24:0] addend_x__2_squeezed;
  wire [7:0] a_bexp__4;
  wire [7:0] incremented_sum__1;
  wire [7:0] MAX_EXPONENT;
  wire [22:0] a_fraction__1;
  wire [7:0] b_bexp__5;
  wire [7:0] MAX_EXPONENT__1;
  wire [22:0] b_fraction__5;
  wire p2_data_enable;
  wire p2_not_valid;
  wire [9:0] wide_exponent;
  wire do_round_up;
  wire [24:0] add_21563;
  wire [3:0] leading_zeroes__0_to_4;
  wire nor_21345;
  wire nor_21346;
  wire nor_21348;
  wire nor_21349;
  wire nor_21354;
  wire nor_21355;
  wire nor_21360;
  wire nor_21363;
  wire nor_21364;
  wire nor_21365;
  wire nor_21371;
  wire [7:0] a_bexpbs_difference__2;
  wire eq_21229;
  wire eq_21230;
  wire eq_21231;
  wire eq_21232;
  wire p1_enable;
  wire and_reduce_21626;
  wire [9:0] wide_exponent__1;
  wire [24:0] rounded_fraction_squeezed_portion_3_width_25;
  wire [4:0] leading_zeroes;
  wire nor_21372;
  wire and_21373;
  wire and_21375;
  wire nor_21380;
  wire and_21381;
  wire nor_21384;
  wire and_21388;
  wire nor_21389;
  wire and_21393;
  wire nor_21395;
  wire [25:0] add_21281;
  wire [23:0] fraction_x;
  wire a_sign__1;
  wire b_sign__3;
  wire [7:0] b_bexp__4;
  wire p1_data_enable;
  wire p1_not_valid;
  wire rounding_carry;
  wire [2:0] fraction_shift__2;
  wire [2:0] fraction_shift__4;
  wire [28:0] cancel_fraction;
  wire and_21402;
  wire and_21420;
  wire [23:0] fraction_x__1;
  wire [2:0] addend_x__2_squeezed_const_lsb_bits__1;
  wire [23:0] fraction_y;
  wire [23:0] sign_ext_21201;
  wire [27:0] add_21220;
  wire [7:0] a_bexp__2;
  wire p0_enable;
  wire p0_all_active_inputs_valid;
  wire [27:0] rounded_fraction;
  wire [2:0] fraction_shift__1;
  wire [26:0] cancel_fraction__1;
  wire [26:0] carry_fraction__1;
  wire and_21438;
  wire and_21440;
  wire nor_21446;
  wire and_21447;
  wire [1:0] priority_sel_21454;
  wire [27:0] concat_21286;
  wire fraction_is_zero;
  wire [27:0] wide_x;
  wire [23:0] fraction_y__1;
  wire [2:0] addend_x__2_squeezed_const_lsb_bits;
  wire has_pos_inf;
  wire has_neg_inf;
  wire p0_data_enable;
  wire rhs_valid_inv;
  wire lhs_valid_inv;
  wire [22:0] FRACTION_HIGH_BIT;
  wire [7:0] MAX_EXPONENT__2;
  wire [8:0] add_21571;
  wire [27:0] shrl_21577;
  wire [26:0] shifted_fraction;
  wire result_sign__1;
  wire [27:0] neg_21212;
  wire [27:0] wide_y;
  wire [8:0] sum__1;
  wire b_sign__2;
  wire rhs_valid_load_en;
  wire lhs_valid_load_en;
  wire [22:0] result_fraction__4;
  wire [22:0] result_fraction__3;
  wire [7:0] result_exponent__2;
  wire [8:0] wide_exponent__2;
  wire [9:0] concat_21572;
  wire [22:0] result_fraction;
  wire [2:0] normal_chunk;
  wire [1:0] half_way_chunk;
  wire [23:0] bit_slice_21532;
  wire nor_21473;
  wire and_21474;
  wire [2:0] priority_sel_21475;
  wire [1:0] priority_sel_21476;
  wire [2:0] priority_sel_21477;
  wire or_21478;
  wire result_sign__2;
  wire [27:0] abs_fraction__1;
  wire not_21297;
  wire result_sign;
  wire xor_21216;
  wire [24:0] wide_x_squeezed;
  wire [24:0] bit_slice_21218;
  wire [27:0] shrl_21219;
  wire sticky;
  wire is_operand_inf;
  wire and_21249;
  wire is_result_nan;
  wire not_21251;
  wire bit_slice_21156;
  wire [22:0] b_fraction__4;
  wire [22:0] tuple_index_21158;
  wire [7:0] bit_slice_21159;
  wire not_21161;
  wire tuple_index_21162;
  wire rhs_load_en;
  wire lhs_load_en;
  wire [31:0] sum;
  assign result_valid_inv = ~result_valid_reg;
  assign result_valid_load_en = result_ready | result_valid_inv;
  assign result_load_en = p7_valid & result_valid_load_en;
  assign p8_stage_done = p7_valid & result_load_en;
  assign p8_not_valid = ~p7_valid;
  assign p7_enable = p8_stage_done | p8_not_valid;
  assign p7_data_enable = p7_enable & p6_valid;
  assign p7_not_valid = ~p6_valid;
  assign p6_enable = p7_data_enable | p7_not_valid;
  assign p6_data_enable = p6_enable & p5_valid;
  assign p6_not_valid = ~p5_valid;
  assign p5_enable = p6_data_enable | p6_not_valid;
  assign p5_data_enable = p5_enable & p4_valid;
  assign p5_not_valid = ~p4_valid;
  assign p4_enable = p5_data_enable | p5_not_valid;
  assign p4_data_enable = p4_enable & p3_valid;
  assign p4_not_valid = ~p3_valid;
  assign p3_enable = p4_data_enable | p4_not_valid;
  assign p3_data_enable = p3_enable & p2_valid;
  assign p3_not_valid = ~p2_valid;
  assign fraction_shift__3 = 3'h4;
  assign p2_enable = p3_data_enable | p3_not_valid;
  assign add_21599 = p5_concat_21572 + 10'h001;
  assign concat_21560 = {1'h0, p4_bit_slice_21532};
  assign carry_bit = p2_abs_fraction__1[27];
  assign addend_x__2_squeezed = p1_xor_21216 ? p1_bit_slice_21218 : p1_wide_x_squeezed;
  assign a_bexp__4 = p0_bit_slice_21156 ? p0_a_bexp__2 : p0_b_bexp__4;
  assign incremented_sum__1 = p0_bit_slice_21159 + 8'h01;
  assign MAX_EXPONENT = 8'hff;
  assign a_fraction__1 = p0_bit_slice_21156 ? p0_tuple_index_21158 : p0_b_fraction__4;
  assign b_bexp__5 = p0_bit_slice_21156 ? p0_b_bexp__4 : p0_a_bexp__2;
  assign MAX_EXPONENT__1 = 8'hff;
  assign b_fraction__5 = p0_bit_slice_21156 ? p0_b_fraction__4 : p0_tuple_index_21158;
  assign p2_data_enable = p2_enable & p1_valid;
  assign p2_not_valid = ~p1_valid;
  assign wide_exponent = add_21599 - {5'h00, p5_and_21474, p5_leading_zeroes__0_to_4};
  assign do_round_up = p4_normal_chunk > fraction_shift__3 | p4_half_way_chunk == 2'h3;
  assign add_21563 = concat_21560 + 25'h000_0001;
  assign leading_zeroes__0_to_4 = priority_sel_4b_2way({p3_nor_21473, p3_and_21474}, {p3_and_21440, p3_priority_sel_21475}, {1'h1, p3_nor_21446, p3_priority_sel_21476}, {p3_and_21438, p3_priority_sel_21477});
  assign nor_21345 = ~(p2_abs_fraction__1[11] | p2_abs_fraction__1[10]);
  assign nor_21346 = ~(p2_abs_fraction__1[9] | p2_abs_fraction__1[8]);
  assign nor_21348 = ~(p2_abs_fraction__1[1] | p2_abs_fraction__1[0]);
  assign nor_21349 = ~(p2_abs_fraction__1[3] | p2_abs_fraction__1[2]);
  assign nor_21354 = ~(p2_abs_fraction__1[5] | p2_abs_fraction__1[4]);
  assign nor_21355 = ~(p2_abs_fraction__1[7] | p2_abs_fraction__1[6]);
  assign nor_21360 = ~(p2_abs_fraction__1[17] | p2_abs_fraction__1[16]);
  assign nor_21363 = ~(p2_abs_fraction__1[13] | p2_abs_fraction__1[12]);
  assign nor_21364 = ~(carry_bit | p2_abs_fraction__1[26]);
  assign nor_21365 = ~(p2_abs_fraction__1[25] | p2_abs_fraction__1[24]);
  assign nor_21371 = ~(p2_abs_fraction__1[21] | p2_abs_fraction__1[20]);
  assign a_bexpbs_difference__2 = p0_bit_slice_21156 ? incremented_sum__1 : ~p0_bit_slice_21159;
  assign eq_21229 = a_bexp__4 == MAX_EXPONENT;
  assign eq_21230 = a_fraction__1 == 23'h00_0000;
  assign eq_21231 = b_bexp__5 == MAX_EXPONENT__1;
  assign eq_21232 = b_fraction__5 == 23'h00_0000;
  assign p1_enable = p2_data_enable | p2_not_valid;
  assign and_reduce_21626 = &p6_wide_exponent__2[7:0];
  assign wide_exponent__1 = wide_exponent & {10{p5_not_21297}};
  assign rounded_fraction_squeezed_portion_3_width_25 = do_round_up ? add_21563 : concat_21560;
  assign leading_zeroes = {p3_and_21474, leading_zeroes__0_to_4};
  assign nor_21372 = ~(p2_abs_fraction__1[23] | p2_abs_fraction__1[22]);
  assign and_21373 = nor_21345 & nor_21346;
  assign and_21375 = nor_21349 & nor_21348;
  assign nor_21380 = ~(p2_abs_fraction__1[7] | p2_abs_fraction__1[6] | nor_21354);
  assign and_21381 = nor_21355 & nor_21354;
  assign nor_21384 = ~(p2_abs_fraction__1[11] | ~p2_abs_fraction__1[10]);
  assign and_21388 = ~(p2_abs_fraction__1[19] | p2_abs_fraction__1[18]) & nor_21360;
  assign nor_21389 = ~(p2_abs_fraction__1[15] | p2_abs_fraction__1[14]);
  assign and_21393 = nor_21364 & nor_21365;
  assign nor_21395 = ~(carry_bit | ~p2_abs_fraction__1[26]);
  assign add_21281 = {{1{addend_x__2_squeezed[24]}}, addend_x__2_squeezed} + {1'h0, p1_shrl_21219[27:3]};
  assign fraction_x = {1'h1, a_fraction__1};
  assign a_sign__1 = p0_bit_slice_21156 ? p0_tuple_index_21162 : p0_not_21161;
  assign b_sign__3 = p0_bit_slice_21156 ? p0_not_21161 : p0_tuple_index_21162;
  assign b_bexp__4 = rhs_reg[30:23];
  assign p1_data_enable = p1_enable & p0_valid;
  assign p1_not_valid = ~p0_valid;
  assign rounding_carry = rounded_fraction_squeezed_portion_3_width_25[24];
  assign fraction_shift__2 = 3'h3;
  assign fraction_shift__4 = 3'h4;
  assign cancel_fraction = leading_zeroes >= 5'h1d ? 29'h0000_0000 : {1'h0, p3_abs_fraction__1} << leading_zeroes;
  assign and_21402 = nor_21372 & nor_21371;
  assign and_21420 = nor_21389 & nor_21363;
  assign fraction_x__1 = fraction_x & {24{a_bexp__4 != 8'h00}};
  assign addend_x__2_squeezed_const_lsb_bits__1 = 3'h0;
  assign fraction_y = {1'h1, b_fraction__5};
  assign sign_ext_21201 = {24{b_bexp__5 != 8'h00}};
  assign add_21220 = (a_bexpbs_difference__2 >= 8'h1c ? 28'h000_0000 : 28'h000_0001 << a_bexpbs_difference__2) + 28'hfff_ffff;
  assign a_bexp__2 = lhs_reg[30:23];
  assign p0_enable = p1_data_enable | p1_not_valid;
  assign p0_all_active_inputs_valid = rhs_valid_reg & lhs_valid_reg;
  assign rounded_fraction = {rounded_fraction_squeezed_portion_3_width_25, p4_normal_chunk};
  assign fraction_shift__1 = rounding_carry ? fraction_shift__4 : fraction_shift__2;
  assign cancel_fraction__1 = cancel_fraction[27:1];
  assign carry_fraction__1 = {p3_abs_fraction__1[27:2], p3_or_21478};
  assign and_21438 = and_21393 & and_21402;
  assign and_21440 = and_21373 & and_21381;
  assign nor_21446 = ~(~and_21388 | and_21420);
  assign and_21447 = and_21388 & and_21420;
  assign priority_sel_21454 = priority_sel_2b_2way({~(carry_bit | p2_abs_fraction__1[26] | nor_21365), and_21393}, {nor_21395, 1'h0}, {1'h1, ~(p2_abs_fraction__1[25] | ~p2_abs_fraction__1[24])}, {nor_21364, nor_21395});
  assign concat_21286 = {add_21281[24:0], p1_shrl_21219[2:1], p1_shrl_21219[0] | p1_sticky};
  assign fraction_is_zero = add_21281 == 26'h000_0000 & ~(p1_shrl_21219[1] | p1_shrl_21219[2]) & ~(p1_shrl_21219[0] | p1_sticky);
  assign wide_x = {1'h0, fraction_x__1, addend_x__2_squeezed_const_lsb_bits__1};
  assign fraction_y__1 = fraction_y & sign_ext_21201;
  assign addend_x__2_squeezed_const_lsb_bits = 3'h0;
  assign has_pos_inf = ~(~eq_21229 | ~eq_21230 | a_sign__1) | ~(~eq_21231 | ~eq_21232 | b_sign__3);
  assign has_neg_inf = eq_21229 & eq_21230 & a_sign__1 | eq_21231 & eq_21232 & b_sign__3;
  assign p0_data_enable = p0_enable & p0_all_active_inputs_valid;
  assign rhs_valid_inv = ~rhs_valid_reg;
  assign lhs_valid_inv = ~lhs_valid_reg;
  assign FRACTION_HIGH_BIT = 23'h40_0000;
  assign MAX_EXPONENT__2 = 8'hff;
  assign add_21571 = {1'h0, p4_a_bexp__4} + {8'h00, rounding_carry};
  assign shrl_21577 = rounded_fraction >> fraction_shift__1;
  assign shifted_fraction = p3_carry_bit ? carry_fraction__1 : cancel_fraction__1;
  assign result_sign__1 = p2_is_operand_inf ? p2_not_21251 : p2_result_sign;
  assign neg_21212 = -wide_x;
  assign wide_y = {1'h0, fraction_y__1, addend_x__2_squeezed_const_lsb_bits};
  assign sum__1 = {1'h0, a_bexp__2} + {1'h0, ~b_bexp__4};
  assign b_sign__2 = rhs_reg[31:31];
  assign rhs_valid_load_en = p0_data_enable | rhs_valid_inv;
  assign lhs_valid_load_en = p0_data_enable | lhs_valid_inv;
  assign result_fraction__4 = p7_is_result_nan ? FRACTION_HIGH_BIT : p7_result_fraction__3;
  assign result_fraction__3 = p6_result_fraction & {23{~(p6_is_operand_inf | p6_wide_exponent__2[8] | and_reduce_21626 | ~((|p6_wide_exponent__2[8:1]) | p6_wide_exponent__2[0]))}};
  assign result_exponent__2 = p6_is_result_nan | p6_is_operand_inf | p6_wide_exponent__2[8] | and_reduce_21626 ? MAX_EXPONENT__2 : p6_wide_exponent__2[7:0];
  assign wide_exponent__2 = wide_exponent__1[8:0] & {9{~wide_exponent__1[9]}};
  assign concat_21572 = {1'h0, add_21571};
  assign result_fraction = shrl_21577[22:0];
  assign normal_chunk = shifted_fraction[2:0];
  assign half_way_chunk = shifted_fraction[3:2];
  assign bit_slice_21532 = shifted_fraction[26:3];
  assign nor_21473 = ~(~and_21438 | and_21447);
  assign and_21474 = and_21438 & and_21447;
  assign priority_sel_21475 = priority_sel_3b_2way({~(~and_21373 | and_21381), and_21440}, {and_21375, priority_sel_2b_2way({~(p2_abs_fraction__1[3] | p2_abs_fraction__1[2] | nor_21348), and_21375}, 2'h0, {1'h1, ~(p2_abs_fraction__1[1] | ~p2_abs_fraction__1[0])}, {nor_21349, ~(p2_abs_fraction__1[3] | ~p2_abs_fraction__1[2])})}, {1'h1, nor_21380, priority_sel_1b_4way({~(p2_abs_fraction__1[7] | ~p2_abs_fraction__1[6]), nor_21355, nor_21380, and_21381}, 1'h0, ~(p2_abs_fraction__1[5] | ~p2_abs_fraction__1[4]), 1'h0, 1'h1, 1'h0)}, {and_21373, priority_sel_2b_2way({~(p2_abs_fraction__1[11] | p2_abs_fraction__1[10] | nor_21346), and_21373}, {nor_21384, 1'h0}, {1'h1, ~(p2_abs_fraction__1[9] | ~p2_abs_fraction__1[8])}, {nor_21345, nor_21384})});
  assign priority_sel_21476 = priority_sel_2b_4way({~(p2_abs_fraction__1[19] | p2_abs_fraction__1[18] | nor_21360), and_21388, nor_21446, and_21447}, 2'h0, {nor_21389, priority_sel_1b_3way({~(p2_abs_fraction__1[15] | ~p2_abs_fraction__1[14]), nor_21389, ~(p2_abs_fraction__1[15] | p2_abs_fraction__1[14] | nor_21363)}, ~(p2_abs_fraction__1[13] | ~p2_abs_fraction__1[12]), 1'h0, 1'h1, 1'h0)}, 2'h0, {1'h1, ~(p2_abs_fraction__1[17] | ~p2_abs_fraction__1[16])}, {1'h0, ~(p2_abs_fraction__1[19] | ~p2_abs_fraction__1[18])});
  assign priority_sel_21477 = priority_sel_3b_2way({~(~and_21393 | and_21402), and_21438}, {priority_sel_21454, 1'h0}, {1'h1, nor_21372, priority_sel_1b_3way({~(p2_abs_fraction__1[23] | ~p2_abs_fraction__1[22]), nor_21372, ~(p2_abs_fraction__1[23] | p2_abs_fraction__1[22] | nor_21371)}, ~(p2_abs_fraction__1[21] | ~p2_abs_fraction__1[20]), 1'h0, 1'h1, 1'h0)}, {and_21393, priority_sel_21454});
  assign or_21478 = p2_abs_fraction__1[1] | p2_abs_fraction__1[0];
  assign result_sign__2 = ~p2_is_result_nan & result_sign__1;
  assign abs_fraction__1 = add_21281[25] ? -concat_21286 : concat_21286;
  assign not_21297 = ~fraction_is_zero;
  assign result_sign = priority_sel_1b_2way({add_21281[25], fraction_is_zero}, p1_and_21249, ~p1_b_sign__3, p1_b_sign__3);
  assign xor_21216 = a_sign__1 ^ b_sign__3;
  assign wide_x_squeezed = {1'h0, fraction_x__1};
  assign bit_slice_21218 = neg_21212[27:3];
  assign shrl_21219 = a_bexpbs_difference__2 >= 8'h1c ? 28'h000_0000 : wide_y >> a_bexpbs_difference__2;
  assign sticky = (fraction_y & sign_ext_21201 & add_21220[26:3]) != 24'h00_0000;
  assign is_operand_inf = eq_21229 & eq_21230 | eq_21231 & eq_21232;
  assign and_21249 = a_sign__1 & b_sign__3;
  assign is_result_nan = ~(~eq_21229 | eq_21230) | ~(~eq_21231 | eq_21232) | has_pos_inf & has_neg_inf;
  assign not_21251 = ~has_pos_inf;
  assign bit_slice_21156 = sum__1[8];
  assign b_fraction__4 = rhs_reg[22:0];
  assign tuple_index_21158 = lhs_reg[22:0];
  assign bit_slice_21159 = sum__1[7:0];
  assign not_21161 = ~b_sign__2;
  assign tuple_index_21162 = lhs_reg[31:31];
  assign rhs_load_en = rhs_valid & rhs_valid_load_en;
  assign lhs_load_en = lhs_valid & lhs_valid_load_en;
  assign sum = {p7_result_sign__2, p7_result_exponent__2, result_fraction__4};
  always @ (posedge clk) begin
    if (rst) begin
      p0_b_bexp__4 <= 8'h00;
      p0_a_bexp__2 <= 8'h00;
      p0_bit_slice_21156 <= 1'h0;
      p0_b_fraction__4 <= 23'h00_0000;
      p0_tuple_index_21158 <= 23'h00_0000;
      p0_bit_slice_21159 <= 8'h00;
      p0_not_21161 <= 1'h0;
      p0_tuple_index_21162 <= 1'h0;
      p1_a_bexp__4 <= 8'h00;
      p1_b_sign__3 <= 1'h0;
      p1_xor_21216 <= 1'h0;
      p1_wide_x_squeezed <= 25'h000_0000;
      p1_bit_slice_21218 <= 25'h000_0000;
      p1_shrl_21219 <= 28'h000_0000;
      p1_sticky <= 1'h0;
      p1_is_operand_inf <= 1'h0;
      p1_and_21249 <= 1'h0;
      p1_is_result_nan <= 1'h0;
      p1_not_21251 <= 1'h0;
      p2_a_bexp__4 <= 8'h00;
      p2_abs_fraction__1 <= 28'h000_0000;
      p2_not_21297 <= 1'h0;
      p2_is_operand_inf <= 1'h0;
      p2_is_result_nan <= 1'h0;
      p2_result_sign <= 1'h0;
      p2_not_21251 <= 1'h0;
      p3_a_bexp__4 <= 8'h00;
      p3_abs_fraction__1 <= 28'h000_0000;
      p3_carry_bit <= 1'h0;
      p3_and_21438 <= 1'h0;
      p3_and_21440 <= 1'h0;
      p3_nor_21446 <= 1'h0;
      p3_nor_21473 <= 1'h0;
      p3_and_21474 <= 1'h0;
      p3_priority_sel_21475 <= 3'h0;
      p3_priority_sel_21476 <= 2'h0;
      p3_priority_sel_21477 <= 3'h0;
      p3_or_21478 <= 1'h0;
      p3_not_21297 <= 1'h0;
      p3_is_operand_inf <= 1'h0;
      p3_is_result_nan <= 1'h0;
      p3_result_sign__2 <= 1'h0;
      p4_a_bexp__4 <= 8'h00;
      p4_and_21474 <= 1'h0;
      p4_leading_zeroes__0_to_4 <= 4'h0;
      p4_normal_chunk <= 3'h0;
      p4_half_way_chunk <= 2'h0;
      p4_bit_slice_21532 <= 24'h00_0000;
      p4_not_21297 <= 1'h0;
      p4_is_operand_inf <= 1'h0;
      p4_is_result_nan <= 1'h0;
      p4_result_sign__2 <= 1'h0;
      p5_and_21474 <= 1'h0;
      p5_leading_zeroes__0_to_4 <= 4'h0;
      p5_concat_21572 <= 10'h000;
      p5_not_21297 <= 1'h0;
      p5_is_operand_inf <= 1'h0;
      p5_is_result_nan <= 1'h0;
      p5_result_fraction <= 23'h00_0000;
      p5_result_sign__2 <= 1'h0;
      p6_wide_exponent__2 <= 9'h000;
      p6_is_operand_inf <= 1'h0;
      p6_is_result_nan <= 1'h0;
      p6_result_fraction <= 23'h00_0000;
      p6_result_sign__2 <= 1'h0;
      p7_is_result_nan <= 1'h0;
      p7_result_fraction__3 <= 23'h00_0000;
      p7_result_sign__2 <= 1'h0;
      p7_result_exponent__2 <= 8'h00;
      p0_valid <= 1'h0;
      p1_valid <= 1'h0;
      p2_valid <= 1'h0;
      p3_valid <= 1'h0;
      p4_valid <= 1'h0;
      p5_valid <= 1'h0;
      p6_valid <= 1'h0;
      p7_valid <= 1'h0;
      rhs_reg <= rhs_reg_init;
      rhs_valid_reg <= 1'h0;
      lhs_reg <= lhs_reg_init;
      lhs_valid_reg <= 1'h0;
      result_reg <= result_reg_init;
      result_valid_reg <= 1'h0;
    end else begin
      p0_b_bexp__4 <= p0_data_enable ? b_bexp__4 : p0_b_bexp__4;
      p0_a_bexp__2 <= p0_data_enable ? a_bexp__2 : p0_a_bexp__2;
      p0_bit_slice_21156 <= p0_data_enable ? bit_slice_21156 : p0_bit_slice_21156;
      p0_b_fraction__4 <= p0_data_enable ? b_fraction__4 : p0_b_fraction__4;
      p0_tuple_index_21158 <= p0_data_enable ? tuple_index_21158 : p0_tuple_index_21158;
      p0_bit_slice_21159 <= p0_data_enable ? bit_slice_21159 : p0_bit_slice_21159;
      p0_not_21161 <= p0_data_enable ? not_21161 : p0_not_21161;
      p0_tuple_index_21162 <= p0_data_enable ? tuple_index_21162 : p0_tuple_index_21162;
      p1_a_bexp__4 <= p1_data_enable ? a_bexp__4 : p1_a_bexp__4;
      p1_b_sign__3 <= p1_data_enable ? b_sign__3 : p1_b_sign__3;
      p1_xor_21216 <= p1_data_enable ? xor_21216 : p1_xor_21216;
      p1_wide_x_squeezed <= p1_data_enable ? wide_x_squeezed : p1_wide_x_squeezed;
      p1_bit_slice_21218 <= p1_data_enable ? bit_slice_21218 : p1_bit_slice_21218;
      p1_shrl_21219 <= p1_data_enable ? shrl_21219 : p1_shrl_21219;
      p1_sticky <= p1_data_enable ? sticky : p1_sticky;
      p1_is_operand_inf <= p1_data_enable ? is_operand_inf : p1_is_operand_inf;
      p1_and_21249 <= p1_data_enable ? and_21249 : p1_and_21249;
      p1_is_result_nan <= p1_data_enable ? is_result_nan : p1_is_result_nan;
      p1_not_21251 <= p1_data_enable ? not_21251 : p1_not_21251;
      p2_a_bexp__4 <= p2_data_enable ? p1_a_bexp__4 : p2_a_bexp__4;
      p2_abs_fraction__1 <= p2_data_enable ? abs_fraction__1 : p2_abs_fraction__1;
      p2_not_21297 <= p2_data_enable ? not_21297 : p2_not_21297;
      p2_is_operand_inf <= p2_data_enable ? p1_is_operand_inf : p2_is_operand_inf;
      p2_is_result_nan <= p2_data_enable ? p1_is_result_nan : p2_is_result_nan;
      p2_result_sign <= p2_data_enable ? result_sign : p2_result_sign;
      p2_not_21251 <= p2_data_enable ? p1_not_21251 : p2_not_21251;
      p3_a_bexp__4 <= p3_data_enable ? p2_a_bexp__4 : p3_a_bexp__4;
      p3_abs_fraction__1 <= p3_data_enable ? p2_abs_fraction__1 : p3_abs_fraction__1;
      p3_carry_bit <= p3_data_enable ? carry_bit : p3_carry_bit;
      p3_and_21438 <= p3_data_enable ? and_21438 : p3_and_21438;
      p3_and_21440 <= p3_data_enable ? and_21440 : p3_and_21440;
      p3_nor_21446 <= p3_data_enable ? nor_21446 : p3_nor_21446;
      p3_nor_21473 <= p3_data_enable ? nor_21473 : p3_nor_21473;
      p3_and_21474 <= p3_data_enable ? and_21474 : p3_and_21474;
      p3_priority_sel_21475 <= p3_data_enable ? priority_sel_21475 : p3_priority_sel_21475;
      p3_priority_sel_21476 <= p3_data_enable ? priority_sel_21476 : p3_priority_sel_21476;
      p3_priority_sel_21477 <= p3_data_enable ? priority_sel_21477 : p3_priority_sel_21477;
      p3_or_21478 <= p3_data_enable ? or_21478 : p3_or_21478;
      p3_not_21297 <= p3_data_enable ? p2_not_21297 : p3_not_21297;
      p3_is_operand_inf <= p3_data_enable ? p2_is_operand_inf : p3_is_operand_inf;
      p3_is_result_nan <= p3_data_enable ? p2_is_result_nan : p3_is_result_nan;
      p3_result_sign__2 <= p3_data_enable ? result_sign__2 : p3_result_sign__2;
      p4_a_bexp__4 <= p4_data_enable ? p3_a_bexp__4 : p4_a_bexp__4;
      p4_and_21474 <= p4_data_enable ? p3_and_21474 : p4_and_21474;
      p4_leading_zeroes__0_to_4 <= p4_data_enable ? leading_zeroes__0_to_4 : p4_leading_zeroes__0_to_4;
      p4_normal_chunk <= p4_data_enable ? normal_chunk : p4_normal_chunk;
      p4_half_way_chunk <= p4_data_enable ? half_way_chunk : p4_half_way_chunk;
      p4_bit_slice_21532 <= p4_data_enable ? bit_slice_21532 : p4_bit_slice_21532;
      p4_not_21297 <= p4_data_enable ? p3_not_21297 : p4_not_21297;
      p4_is_operand_inf <= p4_data_enable ? p3_is_operand_inf : p4_is_operand_inf;
      p4_is_result_nan <= p4_data_enable ? p3_is_result_nan : p4_is_result_nan;
      p4_result_sign__2 <= p4_data_enable ? p3_result_sign__2 : p4_result_sign__2;
      p5_and_21474 <= p5_data_enable ? p4_and_21474 : p5_and_21474;
      p5_leading_zeroes__0_to_4 <= p5_data_enable ? p4_leading_zeroes__0_to_4 : p5_leading_zeroes__0_to_4;
      p5_concat_21572 <= p5_data_enable ? concat_21572 : p5_concat_21572;
      p5_not_21297 <= p5_data_enable ? p4_not_21297 : p5_not_21297;
      p5_is_operand_inf <= p5_data_enable ? p4_is_operand_inf : p5_is_operand_inf;
      p5_is_result_nan <= p5_data_enable ? p4_is_result_nan : p5_is_result_nan;
      p5_result_fraction <= p5_data_enable ? result_fraction : p5_result_fraction;
      p5_result_sign__2 <= p5_data_enable ? p4_result_sign__2 : p5_result_sign__2;
      p6_wide_exponent__2 <= p6_data_enable ? wide_exponent__2 : p6_wide_exponent__2;
      p6_is_operand_inf <= p6_data_enable ? p5_is_operand_inf : p6_is_operand_inf;
      p6_is_result_nan <= p6_data_enable ? p5_is_result_nan : p6_is_result_nan;
      p6_result_fraction <= p6_data_enable ? p5_result_fraction : p6_result_fraction;
      p6_result_sign__2 <= p6_data_enable ? p5_result_sign__2 : p6_result_sign__2;
      p7_is_result_nan <= p7_data_enable ? p6_is_result_nan : p7_is_result_nan;
      p7_result_fraction__3 <= p7_data_enable ? result_fraction__3 : p7_result_fraction__3;
      p7_result_sign__2 <= p7_data_enable ? p6_result_sign__2 : p7_result_sign__2;
      p7_result_exponent__2 <= p7_data_enable ? result_exponent__2 : p7_result_exponent__2;
      p0_valid <= p0_enable ? p0_all_active_inputs_valid : p0_valid;
      p1_valid <= p1_enable ? p0_valid : p1_valid;
      p2_valid <= p2_enable ? p1_valid : p2_valid;
      p3_valid <= p3_enable ? p2_valid : p3_valid;
      p4_valid <= p4_enable ? p3_valid : p4_valid;
      p5_valid <= p5_enable ? p4_valid : p5_valid;
      p6_valid <= p6_enable ? p5_valid : p6_valid;
      p7_valid <= p7_enable ? p6_valid : p7_valid;
      rhs_reg <= rhs_load_en ? rhs : rhs_reg;
      rhs_valid_reg <= rhs_valid_load_en ? rhs_valid : rhs_valid_reg;
      lhs_reg <= lhs_load_en ? lhs : lhs_reg;
      lhs_valid_reg <= lhs_valid_load_en ? lhs_valid : lhs_valid_reg;
      result_reg <= result_load_en ? sum : result_reg;
      result_valid_reg <= result_valid_load_en ? p7_valid : result_valid_reg;
    end
  end
  assign result = result_reg;
  assign result_valid = result_valid_reg;
  assign rhs_ready = rhs_load_en;
  assign lhs_ready = lhs_load_en;
endmodule
