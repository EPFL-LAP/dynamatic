library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity jacobi_1d_imper is
  port (
    A_loadData : in std_logic_vector(31 downto 0);
    B_loadData : in std_logic_vector(31 downto 0);
    A_start_valid : in std_logic;
    B_start_valid : in std_logic;
    start_valid : in std_logic;
    clk : in std_logic;
    rst : in std_logic;
    A_end_ready : in std_logic;
    B_end_ready : in std_logic;
    end_ready : in std_logic;
    A_start_ready : out std_logic;
    B_start_ready : out std_logic;
    start_ready : out std_logic;
    A_end_valid : out std_logic;
    B_end_valid : out std_logic;
    end_valid : out std_logic;
    A_loadEn : out std_logic;
    A_loadAddr : out std_logic_vector(6 downto 0);
    A_storeEn : out std_logic;
    A_storeAddr : out std_logic_vector(6 downto 0);
    A_storeData : out std_logic_vector(31 downto 0);
    B_loadEn : out std_logic;
    B_loadAddr : out std_logic_vector(6 downto 0);
    B_storeEn : out std_logic;
    B_storeAddr : out std_logic_vector(6 downto 0);
    B_storeData : out std_logic_vector(31 downto 0)
  );
end entity;

architecture behavioral of jacobi_1d_imper is

  signal fork0_outs_0_valid : std_logic;
  signal fork0_outs_0_ready : std_logic;
  signal fork0_outs_1_valid : std_logic;
  signal fork0_outs_1_ready : std_logic;
  signal fork0_outs_2_valid : std_logic;
  signal fork0_outs_2_ready : std_logic;
  signal fork0_outs_3_valid : std_logic;
  signal fork0_outs_3_ready : std_logic;
  signal fork0_outs_4_valid : std_logic;
  signal fork0_outs_4_ready : std_logic;
  signal mem_controller0_stDone_0_valid : std_logic;
  signal mem_controller0_stDone_0_ready : std_logic;
  signal mem_controller0_ldData_0 : std_logic_vector(31 downto 0);
  signal mem_controller0_ldData_0_valid : std_logic;
  signal mem_controller0_ldData_0_ready : std_logic;
  signal mem_controller0_memEnd_valid : std_logic;
  signal mem_controller0_memEnd_ready : std_logic;
  signal mem_controller0_loadEn : std_logic;
  signal mem_controller0_loadAddr : std_logic_vector(6 downto 0);
  signal mem_controller0_storeEn : std_logic;
  signal mem_controller0_storeAddr : std_logic_vector(6 downto 0);
  signal mem_controller0_storeData : std_logic_vector(31 downto 0);
  signal mem_controller1_ldData_0 : std_logic_vector(31 downto 0);
  signal mem_controller1_ldData_0_valid : std_logic;
  signal mem_controller1_ldData_0_ready : std_logic;
  signal mem_controller1_ldData_1 : std_logic_vector(31 downto 0);
  signal mem_controller1_ldData_1_valid : std_logic;
  signal mem_controller1_ldData_1_ready : std_logic;
  signal mem_controller1_ldData_2 : std_logic_vector(31 downto 0);
  signal mem_controller1_ldData_2_valid : std_logic;
  signal mem_controller1_ldData_2_ready : std_logic;
  signal mem_controller1_stDone_0_valid : std_logic;
  signal mem_controller1_stDone_0_ready : std_logic;
  signal mem_controller1_memEnd_valid : std_logic;
  signal mem_controller1_memEnd_ready : std_logic;
  signal mem_controller1_loadEn : std_logic;
  signal mem_controller1_loadAddr : std_logic_vector(6 downto 0);
  signal mem_controller1_storeEn : std_logic;
  signal mem_controller1_storeAddr : std_logic_vector(6 downto 0);
  signal mem_controller1_storeData : std_logic_vector(31 downto 0);
  signal constant1_outs : std_logic_vector(10 downto 0);
  signal constant1_outs_valid : std_logic;
  signal constant1_outs_ready : std_logic;
  signal fork1_outs_0 : std_logic_vector(10 downto 0);
  signal fork1_outs_0_valid : std_logic;
  signal fork1_outs_0_ready : std_logic;
  signal fork1_outs_1 : std_logic_vector(10 downto 0);
  signal fork1_outs_1_valid : std_logic;
  signal fork1_outs_1_ready : std_logic;
  signal fork1_outs_2 : std_logic_vector(10 downto 0);
  signal fork1_outs_2_valid : std_logic;
  signal fork1_outs_2_ready : std_logic;
  signal fork1_outs_3 : std_logic_vector(10 downto 0);
  signal fork1_outs_3_valid : std_logic;
  signal fork1_outs_3_ready : std_logic;
  signal fork1_outs_4 : std_logic_vector(10 downto 0);
  signal fork1_outs_4_valid : std_logic;
  signal fork1_outs_4_ready : std_logic;
  signal fork1_outs_5 : std_logic_vector(10 downto 0);
  signal fork1_outs_5_valid : std_logic;
  signal fork1_outs_5_ready : std_logic;
  signal fork1_outs_6 : std_logic_vector(10 downto 0);
  signal fork1_outs_6_valid : std_logic;
  signal fork1_outs_6_ready : std_logic;
  signal fork1_outs_7 : std_logic_vector(10 downto 0);
  signal fork1_outs_7_valid : std_logic;
  signal fork1_outs_7_ready : std_logic;
  signal extsi0_outs : std_logic_vector(31 downto 0);
  signal extsi0_outs_valid : std_logic;
  signal extsi0_outs_ready : std_logic;
  signal extsi1_outs : std_logic_vector(31 downto 0);
  signal extsi1_outs_valid : std_logic;
  signal extsi1_outs_ready : std_logic;
  signal extsi5_outs : std_logic_vector(31 downto 0);
  signal extsi5_outs_valid : std_logic;
  signal extsi5_outs_ready : std_logic;
  signal extsi6_outs : std_logic_vector(31 downto 0);
  signal extsi6_outs_valid : std_logic;
  signal extsi6_outs_ready : std_logic;
  signal constant2_outs : std_logic_vector(0 downto 0);
  signal constant2_outs_valid : std_logic;
  signal constant2_outs_ready : std_logic;
  signal extsi21_outs : std_logic_vector(2 downto 0);
  signal extsi21_outs_valid : std_logic;
  signal extsi21_outs_ready : std_logic;
  signal mux6_outs : std_logic_vector(31 downto 0);
  signal mux6_outs_valid : std_logic;
  signal mux6_outs_ready : std_logic;
  signal mux7_outs : std_logic_vector(31 downto 0);
  signal mux7_outs_valid : std_logic;
  signal mux7_outs_ready : std_logic;
  signal mux9_outs : std_logic_vector(10 downto 0);
  signal mux9_outs_valid : std_logic;
  signal mux9_outs_ready : std_logic;
  signal mux10_outs : std_logic_vector(10 downto 0);
  signal mux10_outs_valid : std_logic;
  signal mux10_outs_ready : std_logic;
  signal mux19_outs : std_logic_vector(10 downto 0);
  signal mux19_outs_valid : std_logic;
  signal mux19_outs_ready : std_logic;
  signal mux21_outs : std_logic_vector(31 downto 0);
  signal mux21_outs_valid : std_logic;
  signal mux21_outs_ready : std_logic;
  signal mux23_outs : std_logic_vector(31 downto 0);
  signal mux23_outs_valid : std_logic;
  signal mux23_outs_ready : std_logic;
  signal mux28_outs : std_logic_vector(10 downto 0);
  signal mux28_outs_valid : std_logic;
  signal mux28_outs_ready : std_logic;
  signal mux37_outs_valid : std_logic;
  signal mux37_outs_ready : std_logic;
  signal init0_outs : std_logic_vector(0 downto 0);
  signal init0_outs_valid : std_logic;
  signal init0_outs_ready : std_logic;
  signal fork2_outs_0 : std_logic_vector(0 downto 0);
  signal fork2_outs_0_valid : std_logic;
  signal fork2_outs_0_ready : std_logic;
  signal fork2_outs_1 : std_logic_vector(0 downto 0);
  signal fork2_outs_1_valid : std_logic;
  signal fork2_outs_1_ready : std_logic;
  signal fork2_outs_2 : std_logic_vector(0 downto 0);
  signal fork2_outs_2_valid : std_logic;
  signal fork2_outs_2_ready : std_logic;
  signal fork2_outs_3 : std_logic_vector(0 downto 0);
  signal fork2_outs_3_valid : std_logic;
  signal fork2_outs_3_ready : std_logic;
  signal fork2_outs_4 : std_logic_vector(0 downto 0);
  signal fork2_outs_4_valid : std_logic;
  signal fork2_outs_4_ready : std_logic;
  signal fork2_outs_5 : std_logic_vector(0 downto 0);
  signal fork2_outs_5_valid : std_logic;
  signal fork2_outs_5_ready : std_logic;
  signal fork2_outs_6 : std_logic_vector(0 downto 0);
  signal fork2_outs_6_valid : std_logic;
  signal fork2_outs_6_ready : std_logic;
  signal fork2_outs_7 : std_logic_vector(0 downto 0);
  signal fork2_outs_7_valid : std_logic;
  signal fork2_outs_7_ready : std_logic;
  signal fork2_outs_8 : std_logic_vector(0 downto 0);
  signal fork2_outs_8_valid : std_logic;
  signal fork2_outs_8_ready : std_logic;
  signal mux0_outs : std_logic_vector(2 downto 0);
  signal mux0_outs_valid : std_logic;
  signal mux0_outs_ready : std_logic;
  signal control_merge0_outs_valid : std_logic;
  signal control_merge0_outs_ready : std_logic;
  signal control_merge0_index : std_logic_vector(0 downto 0);
  signal control_merge0_index_valid : std_logic;
  signal control_merge0_index_ready : std_logic;
  signal fork3_outs_0_valid : std_logic;
  signal fork3_outs_0_ready : std_logic;
  signal fork3_outs_1_valid : std_logic;
  signal fork3_outs_1_ready : std_logic;
  signal constant5_outs : std_logic_vector(1 downto 0);
  signal constant5_outs_valid : std_logic;
  signal constant5_outs_ready : std_logic;
  signal extsi20_outs : std_logic_vector(7 downto 0);
  signal extsi20_outs_valid : std_logic;
  signal extsi20_outs_ready : std_logic;
  signal buffer13_outs : std_logic_vector(2 downto 0);
  signal buffer13_outs_valid : std_logic;
  signal buffer13_outs_ready : std_logic;
  signal cond_br205_trueOut : std_logic_vector(31 downto 0);
  signal cond_br205_trueOut_valid : std_logic;
  signal cond_br205_trueOut_ready : std_logic;
  signal cond_br205_falseOut : std_logic_vector(31 downto 0);
  signal cond_br205_falseOut_valid : std_logic;
  signal cond_br205_falseOut_ready : std_logic;
  signal cond_br206_trueOut_valid : std_logic;
  signal cond_br206_trueOut_ready : std_logic;
  signal cond_br206_falseOut_valid : std_logic;
  signal cond_br206_falseOut_ready : std_logic;
  signal cond_br207_trueOut : std_logic_vector(31 downto 0);
  signal cond_br207_trueOut_valid : std_logic;
  signal cond_br207_trueOut_ready : std_logic;
  signal cond_br207_falseOut : std_logic_vector(31 downto 0);
  signal cond_br207_falseOut_valid : std_logic;
  signal cond_br207_falseOut_ready : std_logic;
  signal buffer37_outs : std_logic_vector(31 downto 0);
  signal buffer37_outs_valid : std_logic;
  signal buffer37_outs_ready : std_logic;
  signal cond_br208_trueOut_valid : std_logic;
  signal cond_br208_trueOut_ready : std_logic;
  signal cond_br208_falseOut_valid : std_logic;
  signal cond_br208_falseOut_ready : std_logic;
  signal buffer38_outs : std_logic_vector(0 downto 0);
  signal buffer38_outs_valid : std_logic;
  signal buffer38_outs_ready : std_logic;
  signal cond_br209_trueOut : std_logic_vector(10 downto 0);
  signal cond_br209_trueOut_valid : std_logic;
  signal cond_br209_trueOut_ready : std_logic;
  signal cond_br209_falseOut : std_logic_vector(10 downto 0);
  signal cond_br209_falseOut_valid : std_logic;
  signal cond_br209_falseOut_ready : std_logic;
  signal cond_br210_trueOut_valid : std_logic;
  signal cond_br210_trueOut_ready : std_logic;
  signal cond_br210_falseOut_valid : std_logic;
  signal cond_br210_falseOut_ready : std_logic;
  signal cond_br211_trueOut : std_logic_vector(31 downto 0);
  signal cond_br211_trueOut_valid : std_logic;
  signal cond_br211_trueOut_ready : std_logic;
  signal cond_br211_falseOut : std_logic_vector(31 downto 0);
  signal cond_br211_falseOut_valid : std_logic;
  signal cond_br211_falseOut_ready : std_logic;
  signal cond_br212_trueOut : std_logic_vector(7 downto 0);
  signal cond_br212_trueOut_valid : std_logic;
  signal cond_br212_trueOut_ready : std_logic;
  signal cond_br212_falseOut : std_logic_vector(7 downto 0);
  signal cond_br212_falseOut_valid : std_logic;
  signal cond_br212_falseOut_ready : std_logic;
  signal cond_br213_trueOut : std_logic_vector(31 downto 0);
  signal cond_br213_trueOut_valid : std_logic;
  signal cond_br213_trueOut_ready : std_logic;
  signal cond_br213_falseOut : std_logic_vector(31 downto 0);
  signal cond_br213_falseOut_valid : std_logic;
  signal cond_br213_falseOut_ready : std_logic;
  signal cond_br214_trueOut_valid : std_logic;
  signal cond_br214_trueOut_ready : std_logic;
  signal cond_br214_falseOut_valid : std_logic;
  signal cond_br214_falseOut_ready : std_logic;
  signal cond_br215_trueOut_valid : std_logic;
  signal cond_br215_trueOut_ready : std_logic;
  signal cond_br215_falseOut_valid : std_logic;
  signal cond_br215_falseOut_ready : std_logic;
  signal cond_br216_trueOut_valid : std_logic;
  signal cond_br216_trueOut_ready : std_logic;
  signal cond_br216_falseOut_valid : std_logic;
  signal cond_br216_falseOut_ready : std_logic;
  signal cond_br217_trueOut : std_logic_vector(31 downto 0);
  signal cond_br217_trueOut_valid : std_logic;
  signal cond_br217_trueOut_ready : std_logic;
  signal cond_br217_falseOut : std_logic_vector(31 downto 0);
  signal cond_br217_falseOut_valid : std_logic;
  signal cond_br217_falseOut_ready : std_logic;
  signal cond_br218_trueOut : std_logic_vector(10 downto 0);
  signal cond_br218_trueOut_valid : std_logic;
  signal cond_br218_trueOut_ready : std_logic;
  signal cond_br218_falseOut : std_logic_vector(10 downto 0);
  signal cond_br218_falseOut_valid : std_logic;
  signal cond_br218_falseOut_ready : std_logic;
  signal cond_br219_trueOut_valid : std_logic;
  signal cond_br219_trueOut_ready : std_logic;
  signal cond_br219_falseOut_valid : std_logic;
  signal cond_br219_falseOut_ready : std_logic;
  signal cond_br220_trueOut : std_logic_vector(8 downto 0);
  signal cond_br220_trueOut_valid : std_logic;
  signal cond_br220_trueOut_ready : std_logic;
  signal cond_br220_falseOut : std_logic_vector(8 downto 0);
  signal cond_br220_falseOut_valid : std_logic;
  signal cond_br220_falseOut_ready : std_logic;
  signal cond_br221_trueOut_valid : std_logic;
  signal cond_br221_trueOut_ready : std_logic;
  signal cond_br221_falseOut_valid : std_logic;
  signal cond_br221_falseOut_ready : std_logic;
  signal buffer57_outs : std_logic_vector(0 downto 0);
  signal buffer57_outs_valid : std_logic;
  signal buffer57_outs_ready : std_logic;
  signal cond_br222_trueOut : std_logic_vector(10 downto 0);
  signal cond_br222_trueOut_valid : std_logic;
  signal cond_br222_trueOut_ready : std_logic;
  signal cond_br222_falseOut : std_logic_vector(10 downto 0);
  signal cond_br222_falseOut_valid : std_logic;
  signal cond_br222_falseOut_ready : std_logic;
  signal cond_br223_trueOut_valid : std_logic;
  signal cond_br223_trueOut_ready : std_logic;
  signal cond_br223_falseOut_valid : std_logic;
  signal cond_br223_falseOut_ready : std_logic;
  signal cond_br224_trueOut : std_logic_vector(31 downto 0);
  signal cond_br224_trueOut_valid : std_logic;
  signal cond_br224_trueOut_ready : std_logic;
  signal cond_br224_falseOut : std_logic_vector(31 downto 0);
  signal cond_br224_falseOut_valid : std_logic;
  signal cond_br224_falseOut_ready : std_logic;
  signal cond_br225_trueOut : std_logic_vector(31 downto 0);
  signal cond_br225_trueOut_valid : std_logic;
  signal cond_br225_trueOut_ready : std_logic;
  signal cond_br225_falseOut : std_logic_vector(31 downto 0);
  signal cond_br225_falseOut_valid : std_logic;
  signal cond_br225_falseOut_ready : std_logic;
  signal cond_br226_trueOut_valid : std_logic;
  signal cond_br226_trueOut_ready : std_logic;
  signal cond_br226_falseOut_valid : std_logic;
  signal cond_br226_falseOut_ready : std_logic;
  signal cond_br227_trueOut : std_logic_vector(31 downto 0);
  signal cond_br227_trueOut_valid : std_logic;
  signal cond_br227_trueOut_ready : std_logic;
  signal cond_br227_falseOut : std_logic_vector(31 downto 0);
  signal cond_br227_falseOut_valid : std_logic;
  signal cond_br227_falseOut_ready : std_logic;
  signal cond_br228_trueOut_valid : std_logic;
  signal cond_br228_trueOut_ready : std_logic;
  signal cond_br228_falseOut_valid : std_logic;
  signal cond_br228_falseOut_ready : std_logic;
  signal cond_br229_trueOut_valid : std_logic;
  signal cond_br229_trueOut_ready : std_logic;
  signal cond_br229_falseOut_valid : std_logic;
  signal cond_br229_falseOut_ready : std_logic;
  signal buffer66_outs : std_logic_vector(0 downto 0);
  signal buffer66_outs_valid : std_logic;
  signal buffer66_outs_ready : std_logic;
  signal cond_br230_trueOut : std_logic_vector(7 downto 0);
  signal cond_br230_trueOut_valid : std_logic;
  signal cond_br230_trueOut_ready : std_logic;
  signal cond_br230_falseOut : std_logic_vector(7 downto 0);
  signal cond_br230_falseOut_valid : std_logic;
  signal cond_br230_falseOut_ready : std_logic;
  signal buffer68_outs : std_logic_vector(7 downto 0);
  signal buffer68_outs_valid : std_logic;
  signal buffer68_outs_ready : std_logic;
  signal cond_br231_trueOut_valid : std_logic;
  signal cond_br231_trueOut_ready : std_logic;
  signal cond_br231_falseOut_valid : std_logic;
  signal cond_br231_falseOut_ready : std_logic;
  signal cond_br232_trueOut : std_logic_vector(31 downto 0);
  signal cond_br232_trueOut_valid : std_logic;
  signal cond_br232_trueOut_ready : std_logic;
  signal cond_br232_falseOut : std_logic_vector(31 downto 0);
  signal cond_br232_falseOut_valid : std_logic;
  signal cond_br232_falseOut_ready : std_logic;
  signal cond_br233_trueOut : std_logic_vector(10 downto 0);
  signal cond_br233_trueOut_valid : std_logic;
  signal cond_br233_trueOut_ready : std_logic;
  signal cond_br233_falseOut : std_logic_vector(10 downto 0);
  signal cond_br233_falseOut_valid : std_logic;
  signal cond_br233_falseOut_ready : std_logic;
  signal init40_outs : std_logic_vector(0 downto 0);
  signal init40_outs_valid : std_logic;
  signal init40_outs_ready : std_logic;
  signal fork4_outs_0 : std_logic_vector(0 downto 0);
  signal fork4_outs_0_valid : std_logic;
  signal fork4_outs_0_ready : std_logic;
  signal fork4_outs_1 : std_logic_vector(0 downto 0);
  signal fork4_outs_1_valid : std_logic;
  signal fork4_outs_1_ready : std_logic;
  signal fork4_outs_2 : std_logic_vector(0 downto 0);
  signal fork4_outs_2_valid : std_logic;
  signal fork4_outs_2_ready : std_logic;
  signal fork4_outs_3 : std_logic_vector(0 downto 0);
  signal fork4_outs_3_valid : std_logic;
  signal fork4_outs_3_ready : std_logic;
  signal fork4_outs_4 : std_logic_vector(0 downto 0);
  signal fork4_outs_4_valid : std_logic;
  signal fork4_outs_4_ready : std_logic;
  signal fork4_outs_5 : std_logic_vector(0 downto 0);
  signal fork4_outs_5_valid : std_logic;
  signal fork4_outs_5_ready : std_logic;
  signal fork4_outs_6 : std_logic_vector(0 downto 0);
  signal fork4_outs_6_valid : std_logic;
  signal fork4_outs_6_ready : std_logic;
  signal fork4_outs_7 : std_logic_vector(0 downto 0);
  signal fork4_outs_7_valid : std_logic;
  signal fork4_outs_7_ready : std_logic;
  signal fork4_outs_8 : std_logic_vector(0 downto 0);
  signal fork4_outs_8_valid : std_logic;
  signal fork4_outs_8_ready : std_logic;
  signal buffer12_outs_valid : std_logic;
  signal buffer12_outs_ready : std_logic;
  signal mux45_outs_valid : std_logic;
  signal mux45_outs_ready : std_logic;
  signal buffer14_outs_valid : std_logic;
  signal buffer14_outs_ready : std_logic;
  signal buffer15_outs_valid : std_logic;
  signal buffer15_outs_ready : std_logic;
  signal fork5_outs_0_valid : std_logic;
  signal fork5_outs_0_ready : std_logic;
  signal fork5_outs_1_valid : std_logic;
  signal fork5_outs_1_ready : std_logic;
  signal fork5_outs_2_valid : std_logic;
  signal fork5_outs_2_ready : std_logic;
  signal fork5_outs_3_valid : std_logic;
  signal fork5_outs_3_ready : std_logic;
  signal fork5_outs_4_valid : std_logic;
  signal fork5_outs_4_ready : std_logic;
  signal fork5_outs_5_valid : std_logic;
  signal fork5_outs_5_ready : std_logic;
  signal fork5_outs_6_valid : std_logic;
  signal fork5_outs_6_ready : std_logic;
  signal fork5_outs_7_valid : std_logic;
  signal fork5_outs_7_ready : std_logic;
  signal fork5_outs_8_valid : std_logic;
  signal fork5_outs_8_ready : std_logic;
  signal fork5_outs_9_valid : std_logic;
  signal fork5_outs_9_ready : std_logic;
  signal fork5_outs_10_valid : std_logic;
  signal fork5_outs_10_ready : std_logic;
  signal fork5_outs_11_valid : std_logic;
  signal fork5_outs_11_ready : std_logic;
  signal fork5_outs_12_valid : std_logic;
  signal fork5_outs_12_ready : std_logic;
  signal mux48_outs : std_logic_vector(31 downto 0);
  signal mux48_outs_valid : std_logic;
  signal mux48_outs_ready : std_logic;
  signal buffer16_outs : std_logic_vector(31 downto 0);
  signal buffer16_outs_valid : std_logic;
  signal buffer16_outs_ready : std_logic;
  signal buffer17_outs : std_logic_vector(31 downto 0);
  signal buffer17_outs_valid : std_logic;
  signal buffer17_outs_ready : std_logic;
  signal fork6_outs_0 : std_logic_vector(31 downto 0);
  signal fork6_outs_0_valid : std_logic;
  signal fork6_outs_0_ready : std_logic;
  signal fork6_outs_1 : std_logic_vector(31 downto 0);
  signal fork6_outs_1_valid : std_logic;
  signal fork6_outs_1_ready : std_logic;
  signal mux51_outs : std_logic_vector(10 downto 0);
  signal mux51_outs_valid : std_logic;
  signal mux51_outs_ready : std_logic;
  signal buffer18_outs : std_logic_vector(10 downto 0);
  signal buffer18_outs_valid : std_logic;
  signal buffer18_outs_ready : std_logic;
  signal buffer19_outs : std_logic_vector(10 downto 0);
  signal buffer19_outs_valid : std_logic;
  signal buffer19_outs_ready : std_logic;
  signal fork7_outs_0 : std_logic_vector(10 downto 0);
  signal fork7_outs_0_valid : std_logic;
  signal fork7_outs_0_ready : std_logic;
  signal fork7_outs_1 : std_logic_vector(10 downto 0);
  signal fork7_outs_1_valid : std_logic;
  signal fork7_outs_1_ready : std_logic;
  signal extsi22_outs : std_logic_vector(31 downto 0);
  signal extsi22_outs_valid : std_logic;
  signal extsi22_outs_ready : std_logic;
  signal mux52_outs : std_logic_vector(10 downto 0);
  signal mux52_outs_valid : std_logic;
  signal mux52_outs_ready : std_logic;
  signal buffer20_outs : std_logic_vector(10 downto 0);
  signal buffer20_outs_valid : std_logic;
  signal buffer20_outs_ready : std_logic;
  signal buffer21_outs : std_logic_vector(10 downto 0);
  signal buffer21_outs_valid : std_logic;
  signal buffer21_outs_ready : std_logic;
  signal fork8_outs_0 : std_logic_vector(10 downto 0);
  signal fork8_outs_0_valid : std_logic;
  signal fork8_outs_0_ready : std_logic;
  signal fork8_outs_1 : std_logic_vector(10 downto 0);
  signal fork8_outs_1_valid : std_logic;
  signal fork8_outs_1_ready : std_logic;
  signal extsi23_outs : std_logic_vector(31 downto 0);
  signal extsi23_outs_valid : std_logic;
  signal extsi23_outs_ready : std_logic;
  signal mux54_outs : std_logic_vector(31 downto 0);
  signal mux54_outs_valid : std_logic;
  signal mux54_outs_ready : std_logic;
  signal buffer22_outs : std_logic_vector(31 downto 0);
  signal buffer22_outs_valid : std_logic;
  signal buffer22_outs_ready : std_logic;
  signal buffer23_outs : std_logic_vector(31 downto 0);
  signal buffer23_outs_valid : std_logic;
  signal buffer23_outs_ready : std_logic;
  signal fork9_outs_0 : std_logic_vector(31 downto 0);
  signal fork9_outs_0_valid : std_logic;
  signal fork9_outs_0_ready : std_logic;
  signal fork9_outs_1 : std_logic_vector(31 downto 0);
  signal fork9_outs_1_valid : std_logic;
  signal fork9_outs_1_ready : std_logic;
  signal mux56_outs : std_logic_vector(31 downto 0);
  signal mux56_outs_valid : std_logic;
  signal mux56_outs_ready : std_logic;
  signal buffer24_outs : std_logic_vector(31 downto 0);
  signal buffer24_outs_valid : std_logic;
  signal buffer24_outs_ready : std_logic;
  signal buffer25_outs : std_logic_vector(31 downto 0);
  signal buffer25_outs_valid : std_logic;
  signal buffer25_outs_ready : std_logic;
  signal fork10_outs_0 : std_logic_vector(31 downto 0);
  signal fork10_outs_0_valid : std_logic;
  signal fork10_outs_0_ready : std_logic;
  signal fork10_outs_1 : std_logic_vector(31 downto 0);
  signal fork10_outs_1_valid : std_logic;
  signal fork10_outs_1_ready : std_logic;
  signal mux57_outs : std_logic_vector(31 downto 0);
  signal mux57_outs_valid : std_logic;
  signal mux57_outs_ready : std_logic;
  signal buffer26_outs : std_logic_vector(31 downto 0);
  signal buffer26_outs_valid : std_logic;
  signal buffer26_outs_ready : std_logic;
  signal buffer27_outs : std_logic_vector(31 downto 0);
  signal buffer27_outs_valid : std_logic;
  signal buffer27_outs_ready : std_logic;
  signal fork11_outs_0 : std_logic_vector(31 downto 0);
  signal fork11_outs_0_valid : std_logic;
  signal fork11_outs_0_ready : std_logic;
  signal fork11_outs_1 : std_logic_vector(31 downto 0);
  signal fork11_outs_1_valid : std_logic;
  signal fork11_outs_1_ready : std_logic;
  signal mux58_outs : std_logic_vector(10 downto 0);
  signal mux58_outs_valid : std_logic;
  signal mux58_outs_ready : std_logic;
  signal buffer28_outs : std_logic_vector(10 downto 0);
  signal buffer28_outs_valid : std_logic;
  signal buffer28_outs_ready : std_logic;
  signal buffer29_outs : std_logic_vector(10 downto 0);
  signal buffer29_outs_valid : std_logic;
  signal buffer29_outs_ready : std_logic;
  signal fork12_outs_0 : std_logic_vector(10 downto 0);
  signal fork12_outs_0_valid : std_logic;
  signal fork12_outs_0_ready : std_logic;
  signal fork12_outs_1 : std_logic_vector(10 downto 0);
  signal fork12_outs_1_valid : std_logic;
  signal fork12_outs_1_ready : std_logic;
  signal extsi24_outs : std_logic_vector(31 downto 0);
  signal extsi24_outs_valid : std_logic;
  signal extsi24_outs_ready : std_logic;
  signal mux60_outs : std_logic_vector(10 downto 0);
  signal mux60_outs_valid : std_logic;
  signal mux60_outs_ready : std_logic;
  signal buffer30_outs : std_logic_vector(10 downto 0);
  signal buffer30_outs_valid : std_logic;
  signal buffer30_outs_ready : std_logic;
  signal buffer31_outs : std_logic_vector(10 downto 0);
  signal buffer31_outs_valid : std_logic;
  signal buffer31_outs_ready : std_logic;
  signal fork13_outs_0 : std_logic_vector(10 downto 0);
  signal fork13_outs_0_valid : std_logic;
  signal fork13_outs_0_ready : std_logic;
  signal fork13_outs_1 : std_logic_vector(10 downto 0);
  signal fork13_outs_1_valid : std_logic;
  signal fork13_outs_1_ready : std_logic;
  signal extsi25_outs : std_logic_vector(31 downto 0);
  signal extsi25_outs_valid : std_logic;
  signal extsi25_outs_ready : std_logic;
  signal unbundle3_outs_0_valid : std_logic;
  signal unbundle3_outs_0_ready : std_logic;
  signal unbundle3_outs_1 : std_logic_vector(31 downto 0);
  signal unbundle4_outs_0_valid : std_logic;
  signal unbundle4_outs_0_ready : std_logic;
  signal unbundle4_outs_1 : std_logic_vector(31 downto 0);
  signal unbundle5_outs_0_valid : std_logic;
  signal unbundle5_outs_0_ready : std_logic;
  signal unbundle5_outs_1 : std_logic_vector(31 downto 0);
  signal mux1_outs : std_logic_vector(7 downto 0);
  signal mux1_outs_valid : std_logic;
  signal mux1_outs_ready : std_logic;
  signal buffer32_outs : std_logic_vector(7 downto 0);
  signal buffer32_outs_valid : std_logic;
  signal buffer32_outs_ready : std_logic;
  signal buffer33_outs : std_logic_vector(7 downto 0);
  signal buffer33_outs_valid : std_logic;
  signal buffer33_outs_ready : std_logic;
  signal fork14_outs_0 : std_logic_vector(7 downto 0);
  signal fork14_outs_0_valid : std_logic;
  signal fork14_outs_0_ready : std_logic;
  signal fork14_outs_1 : std_logic_vector(7 downto 0);
  signal fork14_outs_1_valid : std_logic;
  signal fork14_outs_1_ready : std_logic;
  signal fork14_outs_2 : std_logic_vector(7 downto 0);
  signal fork14_outs_2_valid : std_logic;
  signal fork14_outs_2_ready : std_logic;
  signal fork14_outs_3 : std_logic_vector(7 downto 0);
  signal fork14_outs_3_valid : std_logic;
  signal fork14_outs_3_ready : std_logic;
  signal fork14_outs_4 : std_logic_vector(7 downto 0);
  signal fork14_outs_4_valid : std_logic;
  signal fork14_outs_4_ready : std_logic;
  signal extsi26_outs : std_logic_vector(8 downto 0);
  signal extsi26_outs_valid : std_logic;
  signal extsi26_outs_ready : std_logic;
  signal extsi27_outs : std_logic_vector(8 downto 0);
  signal extsi27_outs_valid : std_logic;
  signal extsi27_outs_ready : std_logic;
  signal extsi28_outs : std_logic_vector(31 downto 0);
  signal extsi28_outs_valid : std_logic;
  signal extsi28_outs_ready : std_logic;
  signal fork15_outs_0 : std_logic_vector(31 downto 0);
  signal fork15_outs_0_valid : std_logic;
  signal fork15_outs_0_ready : std_logic;
  signal fork15_outs_1 : std_logic_vector(31 downto 0);
  signal fork15_outs_1_valid : std_logic;
  signal fork15_outs_1_ready : std_logic;
  signal fork15_outs_2 : std_logic_vector(31 downto 0);
  signal fork15_outs_2_valid : std_logic;
  signal fork15_outs_2_ready : std_logic;
  signal fork15_outs_3 : std_logic_vector(31 downto 0);
  signal fork15_outs_3_valid : std_logic;
  signal fork15_outs_3_ready : std_logic;
  signal fork15_outs_4 : std_logic_vector(31 downto 0);
  signal fork15_outs_4_valid : std_logic;
  signal fork15_outs_4_ready : std_logic;
  signal mux2_outs : std_logic_vector(2 downto 0);
  signal mux2_outs_valid : std_logic;
  signal mux2_outs_ready : std_logic;
  signal control_merge1_outs_valid : std_logic;
  signal control_merge1_outs_ready : std_logic;
  signal control_merge1_index : std_logic_vector(0 downto 0);
  signal control_merge1_index_valid : std_logic;
  signal control_merge1_index_ready : std_logic;
  signal fork16_outs_0 : std_logic_vector(0 downto 0);
  signal fork16_outs_0_valid : std_logic;
  signal fork16_outs_0_ready : std_logic;
  signal fork16_outs_1 : std_logic_vector(0 downto 0);
  signal fork16_outs_1_valid : std_logic;
  signal fork16_outs_1_ready : std_logic;
  signal buffer36_outs_valid : std_logic;
  signal buffer36_outs_ready : std_logic;
  signal fork17_outs_0_valid : std_logic;
  signal fork17_outs_0_ready : std_logic;
  signal fork17_outs_1_valid : std_logic;
  signal fork17_outs_1_ready : std_logic;
  signal constant16_outs : std_logic_vector(1 downto 0);
  signal constant16_outs_valid : std_logic;
  signal constant16_outs_ready : std_logic;
  signal fork18_outs_0 : std_logic_vector(1 downto 0);
  signal fork18_outs_0_valid : std_logic;
  signal fork18_outs_0_ready : std_logic;
  signal fork18_outs_1 : std_logic_vector(1 downto 0);
  signal fork18_outs_1_valid : std_logic;
  signal fork18_outs_1_ready : std_logic;
  signal fork18_outs_2 : std_logic_vector(1 downto 0);
  signal fork18_outs_2_valid : std_logic;
  signal fork18_outs_2_ready : std_logic;
  signal fork18_outs_3 : std_logic_vector(1 downto 0);
  signal fork18_outs_3_valid : std_logic;
  signal fork18_outs_3_ready : std_logic;
  signal extsi29_outs : std_logic_vector(8 downto 0);
  signal extsi29_outs_valid : std_logic;
  signal extsi29_outs_ready : std_logic;
  signal extsi30_outs : std_logic_vector(8 downto 0);
  signal extsi30_outs_valid : std_logic;
  signal extsi30_outs_ready : std_logic;
  signal extsi11_outs : std_logic_vector(31 downto 0);
  signal extsi11_outs_valid : std_logic;
  signal extsi11_outs_ready : std_logic;
  signal source0_outs_valid : std_logic;
  signal source0_outs_ready : std_logic;
  signal constant7_outs : std_logic_vector(31 downto 0);
  signal constant7_outs_valid : std_logic;
  signal constant7_outs_ready : std_logic;
  signal source1_outs_valid : std_logic;
  signal source1_outs_ready : std_logic;
  signal constant18_outs : std_logic_vector(7 downto 0);
  signal constant18_outs_valid : std_logic;
  signal constant18_outs_ready : std_logic;
  signal extsi31_outs : std_logic_vector(8 downto 0);
  signal extsi31_outs_valid : std_logic;
  signal extsi31_outs_ready : std_logic;
  signal source2_outs_valid : std_logic;
  signal source2_outs_ready : std_logic;
  signal constant19_outs : std_logic_vector(1 downto 0);
  signal constant19_outs_valid : std_logic;
  signal constant19_outs_ready : std_logic;
  signal extsi13_outs : std_logic_vector(31 downto 0);
  signal extsi13_outs_valid : std_logic;
  signal extsi13_outs_ready : std_logic;
  signal addi2_result : std_logic_vector(31 downto 0);
  signal addi2_result_valid : std_logic;
  signal addi2_result_ready : std_logic;
  signal buffer39_outs : std_logic_vector(31 downto 0);
  signal buffer39_outs_valid : std_logic;
  signal buffer39_outs_ready : std_logic;
  signal fork19_outs_0 : std_logic_vector(31 downto 0);
  signal fork19_outs_0_valid : std_logic;
  signal fork19_outs_0_ready : std_logic;
  signal fork19_outs_1 : std_logic_vector(31 downto 0);
  signal fork19_outs_1_valid : std_logic;
  signal fork19_outs_1_ready : std_logic;
  signal fork19_outs_2 : std_logic_vector(31 downto 0);
  signal fork19_outs_2_valid : std_logic;
  signal fork19_outs_2_ready : std_logic;
  signal buffer0_outs : std_logic_vector(31 downto 0);
  signal buffer0_outs_valid : std_logic;
  signal buffer0_outs_ready : std_logic;
  signal fork20_outs_0 : std_logic_vector(31 downto 0);
  signal fork20_outs_0_valid : std_logic;
  signal fork20_outs_0_ready : std_logic;
  signal fork20_outs_1 : std_logic_vector(31 downto 0);
  signal fork20_outs_1_valid : std_logic;
  signal fork20_outs_1_ready : std_logic;
  signal init80_outs : std_logic_vector(31 downto 0);
  signal init80_outs_valid : std_logic;
  signal init80_outs_ready : std_logic;
  signal buffer1_outs_valid : std_logic;
  signal buffer1_outs_ready : std_logic;
  signal fork21_outs_0_valid : std_logic;
  signal fork21_outs_0_ready : std_logic;
  signal fork21_outs_1_valid : std_logic;
  signal fork21_outs_1_ready : std_logic;
  signal init81_outs_valid : std_logic;
  signal init81_outs_ready : std_logic;
  signal fork22_outs_0_valid : std_logic;
  signal fork22_outs_0_ready : std_logic;
  signal fork22_outs_1_valid : std_logic;
  signal fork22_outs_1_ready : std_logic;
  signal init82_outs_valid : std_logic;
  signal init82_outs_ready : std_logic;
  signal gate0_outs : std_logic_vector(31 downto 0);
  signal gate0_outs_valid : std_logic;
  signal gate0_outs_ready : std_logic;
  signal fork23_outs_0 : std_logic_vector(31 downto 0);
  signal fork23_outs_0_valid : std_logic;
  signal fork23_outs_0_ready : std_logic;
  signal fork23_outs_1 : std_logic_vector(31 downto 0);
  signal fork23_outs_1_valid : std_logic;
  signal fork23_outs_1_ready : std_logic;
  signal cmpi3_result : std_logic_vector(0 downto 0);
  signal cmpi3_result_valid : std_logic;
  signal cmpi3_result_ready : std_logic;
  signal fork24_outs_0 : std_logic_vector(0 downto 0);
  signal fork24_outs_0_valid : std_logic;
  signal fork24_outs_0_ready : std_logic;
  signal fork24_outs_1 : std_logic_vector(0 downto 0);
  signal fork24_outs_1_valid : std_logic;
  signal fork24_outs_1_ready : std_logic;
  signal cmpi4_result : std_logic_vector(0 downto 0);
  signal cmpi4_result_valid : std_logic;
  signal cmpi4_result_ready : std_logic;
  signal fork25_outs_0 : std_logic_vector(0 downto 0);
  signal fork25_outs_0_valid : std_logic;
  signal fork25_outs_0_ready : std_logic;
  signal fork25_outs_1 : std_logic_vector(0 downto 0);
  signal fork25_outs_1_valid : std_logic;
  signal fork25_outs_1_ready : std_logic;
  signal cond_br89_trueOut_valid : std_logic;
  signal cond_br89_trueOut_ready : std_logic;
  signal cond_br89_falseOut_valid : std_logic;
  signal cond_br89_falseOut_ready : std_logic;
  signal cond_br90_trueOut_valid : std_logic;
  signal cond_br90_trueOut_ready : std_logic;
  signal cond_br90_falseOut_valid : std_logic;
  signal cond_br90_falseOut_ready : std_logic;
  signal source7_outs_valid : std_logic;
  signal source7_outs_ready : std_logic;
  signal mux85_outs_valid : std_logic;
  signal mux85_outs_ready : std_logic;
  signal source8_outs_valid : std_logic;
  signal source8_outs_ready : std_logic;
  signal mux86_outs_valid : std_logic;
  signal mux86_outs_ready : std_logic;
  signal buffer40_outs_valid : std_logic;
  signal buffer40_outs_ready : std_logic;
  signal buffer41_outs_valid : std_logic;
  signal buffer41_outs_ready : std_logic;
  signal join0_outs_valid : std_logic;
  signal join0_outs_ready : std_logic;
  signal gate1_outs : std_logic_vector(31 downto 0);
  signal gate1_outs_valid : std_logic;
  signal gate1_outs_ready : std_logic;
  signal trunci0_outs : std_logic_vector(6 downto 0);
  signal trunci0_outs_valid : std_logic;
  signal trunci0_outs_ready : std_logic;
  signal load0_addrOut : std_logic_vector(6 downto 0);
  signal load0_addrOut_valid : std_logic;
  signal load0_addrOut_ready : std_logic;
  signal load0_dataOut : std_logic_vector(31 downto 0);
  signal load0_dataOut_valid : std_logic;
  signal load0_dataOut_ready : std_logic;
  signal fork26_outs_0 : std_logic_vector(31 downto 0);
  signal fork26_outs_0_valid : std_logic;
  signal fork26_outs_0_ready : std_logic;
  signal fork26_outs_1 : std_logic_vector(31 downto 0);
  signal fork26_outs_1_valid : std_logic;
  signal fork26_outs_1_ready : std_logic;
  signal buffer2_outs : std_logic_vector(7 downto 0);
  signal buffer2_outs_valid : std_logic;
  signal buffer2_outs_ready : std_logic;
  signal fork27_outs_0 : std_logic_vector(7 downto 0);
  signal fork27_outs_0_valid : std_logic;
  signal fork27_outs_0_ready : std_logic;
  signal fork27_outs_1 : std_logic_vector(7 downto 0);
  signal fork27_outs_1_valid : std_logic;
  signal fork27_outs_1_ready : std_logic;
  signal extsi32_outs : std_logic_vector(31 downto 0);
  signal extsi32_outs_valid : std_logic;
  signal extsi32_outs_ready : std_logic;
  signal init83_outs : std_logic_vector(31 downto 0);
  signal init83_outs_valid : std_logic;
  signal init83_outs_ready : std_logic;
  signal buffer3_outs_valid : std_logic;
  signal buffer3_outs_ready : std_logic;
  signal fork28_outs_0_valid : std_logic;
  signal fork28_outs_0_ready : std_logic;
  signal fork28_outs_1_valid : std_logic;
  signal fork28_outs_1_ready : std_logic;
  signal init84_outs_valid : std_logic;
  signal init84_outs_ready : std_logic;
  signal fork29_outs_0_valid : std_logic;
  signal fork29_outs_0_ready : std_logic;
  signal fork29_outs_1_valid : std_logic;
  signal fork29_outs_1_ready : std_logic;
  signal init85_outs_valid : std_logic;
  signal init85_outs_ready : std_logic;
  signal gate2_outs : std_logic_vector(31 downto 0);
  signal gate2_outs_valid : std_logic;
  signal gate2_outs_ready : std_logic;
  signal fork30_outs_0 : std_logic_vector(31 downto 0);
  signal fork30_outs_0_valid : std_logic;
  signal fork30_outs_0_ready : std_logic;
  signal fork30_outs_1 : std_logic_vector(31 downto 0);
  signal fork30_outs_1_valid : std_logic;
  signal fork30_outs_1_ready : std_logic;
  signal cmpi5_result : std_logic_vector(0 downto 0);
  signal cmpi5_result_valid : std_logic;
  signal cmpi5_result_ready : std_logic;
  signal fork31_outs_0 : std_logic_vector(0 downto 0);
  signal fork31_outs_0_valid : std_logic;
  signal fork31_outs_0_ready : std_logic;
  signal fork31_outs_1 : std_logic_vector(0 downto 0);
  signal fork31_outs_1_valid : std_logic;
  signal fork31_outs_1_ready : std_logic;
  signal cmpi6_result : std_logic_vector(0 downto 0);
  signal cmpi6_result_valid : std_logic;
  signal cmpi6_result_ready : std_logic;
  signal fork32_outs_0 : std_logic_vector(0 downto 0);
  signal fork32_outs_0_valid : std_logic;
  signal fork32_outs_0_ready : std_logic;
  signal fork32_outs_1 : std_logic_vector(0 downto 0);
  signal fork32_outs_1_valid : std_logic;
  signal fork32_outs_1_ready : std_logic;
  signal cond_br91_trueOut_valid : std_logic;
  signal cond_br91_trueOut_ready : std_logic;
  signal cond_br91_falseOut_valid : std_logic;
  signal cond_br91_falseOut_ready : std_logic;
  signal cond_br92_trueOut_valid : std_logic;
  signal cond_br92_trueOut_ready : std_logic;
  signal cond_br92_falseOut_valid : std_logic;
  signal cond_br92_falseOut_ready : std_logic;
  signal source9_outs_valid : std_logic;
  signal source9_outs_ready : std_logic;
  signal mux87_outs_valid : std_logic;
  signal mux87_outs_ready : std_logic;
  signal source10_outs_valid : std_logic;
  signal source10_outs_ready : std_logic;
  signal mux88_outs_valid : std_logic;
  signal mux88_outs_ready : std_logic;
  signal buffer42_outs_valid : std_logic;
  signal buffer42_outs_ready : std_logic;
  signal buffer43_outs_valid : std_logic;
  signal buffer43_outs_ready : std_logic;
  signal join1_outs_valid : std_logic;
  signal join1_outs_ready : std_logic;
  signal gate3_outs : std_logic_vector(31 downto 0);
  signal gate3_outs_valid : std_logic;
  signal gate3_outs_ready : std_logic;
  signal trunci1_outs : std_logic_vector(6 downto 0);
  signal trunci1_outs_valid : std_logic;
  signal trunci1_outs_ready : std_logic;
  signal load1_addrOut : std_logic_vector(6 downto 0);
  signal load1_addrOut_valid : std_logic;
  signal load1_addrOut_ready : std_logic;
  signal load1_dataOut : std_logic_vector(31 downto 0);
  signal load1_dataOut_valid : std_logic;
  signal load1_dataOut_ready : std_logic;
  signal fork33_outs_0 : std_logic_vector(31 downto 0);
  signal fork33_outs_0_valid : std_logic;
  signal fork33_outs_0_ready : std_logic;
  signal fork33_outs_1 : std_logic_vector(31 downto 0);
  signal fork33_outs_1_valid : std_logic;
  signal fork33_outs_1_ready : std_logic;
  signal addi0_result : std_logic_vector(31 downto 0);
  signal addi0_result_valid : std_logic;
  signal addi0_result_ready : std_logic;
  signal addi3_result : std_logic_vector(8 downto 0);
  signal addi3_result_valid : std_logic;
  signal addi3_result_ready : std_logic;
  signal buffer45_outs : std_logic_vector(8 downto 0);
  signal buffer45_outs_valid : std_logic;
  signal buffer45_outs_ready : std_logic;
  signal fork34_outs_0 : std_logic_vector(8 downto 0);
  signal fork34_outs_0_valid : std_logic;
  signal fork34_outs_0_ready : std_logic;
  signal fork34_outs_1 : std_logic_vector(8 downto 0);
  signal fork34_outs_1_valid : std_logic;
  signal fork34_outs_1_ready : std_logic;
  signal extsi33_outs : std_logic_vector(31 downto 0);
  signal extsi33_outs_valid : std_logic;
  signal extsi33_outs_ready : std_logic;
  signal buffer123_outs : std_logic_vector(8 downto 0);
  signal buffer123_outs_valid : std_logic;
  signal buffer123_outs_ready : std_logic;
  signal fork35_outs_0 : std_logic_vector(31 downto 0);
  signal fork35_outs_0_valid : std_logic;
  signal fork35_outs_0_ready : std_logic;
  signal fork35_outs_1 : std_logic_vector(31 downto 0);
  signal fork35_outs_1_valid : std_logic;
  signal fork35_outs_1_ready : std_logic;
  signal buffer4_outs : std_logic_vector(8 downto 0);
  signal buffer4_outs_valid : std_logic;
  signal buffer4_outs_ready : std_logic;
  signal fork36_outs_0 : std_logic_vector(8 downto 0);
  signal fork36_outs_0_valid : std_logic;
  signal fork36_outs_0_ready : std_logic;
  signal fork36_outs_1 : std_logic_vector(8 downto 0);
  signal fork36_outs_1_valid : std_logic;
  signal fork36_outs_1_ready : std_logic;
  signal extsi34_outs : std_logic_vector(31 downto 0);
  signal extsi34_outs_valid : std_logic;
  signal extsi34_outs_ready : std_logic;
  signal init86_outs : std_logic_vector(31 downto 0);
  signal init86_outs_valid : std_logic;
  signal init86_outs_ready : std_logic;
  signal buffer5_outs_valid : std_logic;
  signal buffer5_outs_ready : std_logic;
  signal fork37_outs_0_valid : std_logic;
  signal fork37_outs_0_ready : std_logic;
  signal fork37_outs_1_valid : std_logic;
  signal fork37_outs_1_ready : std_logic;
  signal init87_outs_valid : std_logic;
  signal init87_outs_ready : std_logic;
  signal fork38_outs_0_valid : std_logic;
  signal fork38_outs_0_ready : std_logic;
  signal fork38_outs_1_valid : std_logic;
  signal fork38_outs_1_ready : std_logic;
  signal init88_outs_valid : std_logic;
  signal init88_outs_ready : std_logic;
  signal gate4_outs : std_logic_vector(31 downto 0);
  signal gate4_outs_valid : std_logic;
  signal gate4_outs_ready : std_logic;
  signal fork39_outs_0 : std_logic_vector(31 downto 0);
  signal fork39_outs_0_valid : std_logic;
  signal fork39_outs_0_ready : std_logic;
  signal fork39_outs_1 : std_logic_vector(31 downto 0);
  signal fork39_outs_1_valid : std_logic;
  signal fork39_outs_1_ready : std_logic;
  signal cmpi7_result : std_logic_vector(0 downto 0);
  signal cmpi7_result_valid : std_logic;
  signal cmpi7_result_ready : std_logic;
  signal fork40_outs_0 : std_logic_vector(0 downto 0);
  signal fork40_outs_0_valid : std_logic;
  signal fork40_outs_0_ready : std_logic;
  signal fork40_outs_1 : std_logic_vector(0 downto 0);
  signal fork40_outs_1_valid : std_logic;
  signal fork40_outs_1_ready : std_logic;
  signal cmpi8_result : std_logic_vector(0 downto 0);
  signal cmpi8_result_valid : std_logic;
  signal cmpi8_result_ready : std_logic;
  signal fork41_outs_0 : std_logic_vector(0 downto 0);
  signal fork41_outs_0_valid : std_logic;
  signal fork41_outs_0_ready : std_logic;
  signal fork41_outs_1 : std_logic_vector(0 downto 0);
  signal fork41_outs_1_valid : std_logic;
  signal fork41_outs_1_ready : std_logic;
  signal cond_br93_trueOut_valid : std_logic;
  signal cond_br93_trueOut_ready : std_logic;
  signal cond_br93_falseOut_valid : std_logic;
  signal cond_br93_falseOut_ready : std_logic;
  signal cond_br94_trueOut_valid : std_logic;
  signal cond_br94_trueOut_ready : std_logic;
  signal cond_br94_falseOut_valid : std_logic;
  signal cond_br94_falseOut_ready : std_logic;
  signal source11_outs_valid : std_logic;
  signal source11_outs_ready : std_logic;
  signal mux89_outs_valid : std_logic;
  signal mux89_outs_ready : std_logic;
  signal source12_outs_valid : std_logic;
  signal source12_outs_ready : std_logic;
  signal mux90_outs_valid : std_logic;
  signal mux90_outs_ready : std_logic;
  signal buffer46_outs_valid : std_logic;
  signal buffer46_outs_ready : std_logic;
  signal buffer47_outs_valid : std_logic;
  signal buffer47_outs_ready : std_logic;
  signal join2_outs_valid : std_logic;
  signal join2_outs_ready : std_logic;
  signal gate5_outs : std_logic_vector(31 downto 0);
  signal gate5_outs_valid : std_logic;
  signal gate5_outs_ready : std_logic;
  signal buffer134_outs : std_logic_vector(31 downto 0);
  signal buffer134_outs_valid : std_logic;
  signal buffer134_outs_ready : std_logic;
  signal trunci2_outs : std_logic_vector(6 downto 0);
  signal trunci2_outs_valid : std_logic;
  signal trunci2_outs_ready : std_logic;
  signal load2_addrOut : std_logic_vector(6 downto 0);
  signal load2_addrOut_valid : std_logic;
  signal load2_addrOut_ready : std_logic;
  signal load2_dataOut : std_logic_vector(31 downto 0);
  signal load2_dataOut_valid : std_logic;
  signal load2_dataOut_ready : std_logic;
  signal fork42_outs_0 : std_logic_vector(31 downto 0);
  signal fork42_outs_0_valid : std_logic;
  signal fork42_outs_0_ready : std_logic;
  signal fork42_outs_1 : std_logic_vector(31 downto 0);
  signal fork42_outs_1_valid : std_logic;
  signal fork42_outs_1_ready : std_logic;
  signal buffer44_outs : std_logic_vector(31 downto 0);
  signal buffer44_outs_valid : std_logic;
  signal buffer44_outs_ready : std_logic;
  signal addi1_result : std_logic_vector(31 downto 0);
  signal addi1_result_valid : std_logic;
  signal addi1_result_ready : std_logic;
  signal buffer48_outs : std_logic_vector(31 downto 0);
  signal buffer48_outs_valid : std_logic;
  signal buffer48_outs_ready : std_logic;
  signal fork43_outs_0 : std_logic_vector(31 downto 0);
  signal fork43_outs_0_valid : std_logic;
  signal fork43_outs_0_ready : std_logic;
  signal fork43_outs_1 : std_logic_vector(31 downto 0);
  signal fork43_outs_1_valid : std_logic;
  signal fork43_outs_1_ready : std_logic;
  signal shli0_result : std_logic_vector(31 downto 0);
  signal shli0_result_valid : std_logic;
  signal shli0_result_ready : std_logic;
  signal buffer49_outs : std_logic_vector(31 downto 0);
  signal buffer49_outs_valid : std_logic;
  signal buffer49_outs_ready : std_logic;
  signal addi7_result : std_logic_vector(31 downto 0);
  signal addi7_result_valid : std_logic;
  signal addi7_result_ready : std_logic;
  signal buffer6_outs : std_logic_vector(7 downto 0);
  signal buffer6_outs_valid : std_logic;
  signal buffer6_outs_ready : std_logic;
  signal fork44_outs_0 : std_logic_vector(7 downto 0);
  signal fork44_outs_0_valid : std_logic;
  signal fork44_outs_0_ready : std_logic;
  signal fork44_outs_1 : std_logic_vector(7 downto 0);
  signal fork44_outs_1_valid : std_logic;
  signal fork44_outs_1_ready : std_logic;
  signal extsi35_outs : std_logic_vector(31 downto 0);
  signal extsi35_outs_valid : std_logic;
  signal extsi35_outs_ready : std_logic;
  signal init89_outs : std_logic_vector(31 downto 0);
  signal init89_outs_valid : std_logic;
  signal init89_outs_ready : std_logic;
  signal buffer53_outs_valid : std_logic;
  signal buffer53_outs_ready : std_logic;
  signal buffer7_outs_valid : std_logic;
  signal buffer7_outs_ready : std_logic;
  signal fork45_outs_0_valid : std_logic;
  signal fork45_outs_0_ready : std_logic;
  signal fork45_outs_1_valid : std_logic;
  signal fork45_outs_1_ready : std_logic;
  signal init90_outs_valid : std_logic;
  signal init90_outs_ready : std_logic;
  signal fork46_outs_0_valid : std_logic;
  signal fork46_outs_0_ready : std_logic;
  signal fork46_outs_1_valid : std_logic;
  signal fork46_outs_1_ready : std_logic;
  signal init91_outs_valid : std_logic;
  signal init91_outs_ready : std_logic;
  signal gate6_outs : std_logic_vector(31 downto 0);
  signal gate6_outs_valid : std_logic;
  signal gate6_outs_ready : std_logic;
  signal fork47_outs_0 : std_logic_vector(31 downto 0);
  signal fork47_outs_0_valid : std_logic;
  signal fork47_outs_0_ready : std_logic;
  signal fork47_outs_1 : std_logic_vector(31 downto 0);
  signal fork47_outs_1_valid : std_logic;
  signal fork47_outs_1_ready : std_logic;
  signal cmpi9_result : std_logic_vector(0 downto 0);
  signal cmpi9_result_valid : std_logic;
  signal cmpi9_result_ready : std_logic;
  signal fork48_outs_0 : std_logic_vector(0 downto 0);
  signal fork48_outs_0_valid : std_logic;
  signal fork48_outs_0_ready : std_logic;
  signal fork48_outs_1 : std_logic_vector(0 downto 0);
  signal fork48_outs_1_valid : std_logic;
  signal fork48_outs_1_ready : std_logic;
  signal cmpi10_result : std_logic_vector(0 downto 0);
  signal cmpi10_result_valid : std_logic;
  signal cmpi10_result_ready : std_logic;
  signal fork49_outs_0 : std_logic_vector(0 downto 0);
  signal fork49_outs_0_valid : std_logic;
  signal fork49_outs_0_ready : std_logic;
  signal fork49_outs_1 : std_logic_vector(0 downto 0);
  signal fork49_outs_1_valid : std_logic;
  signal fork49_outs_1_ready : std_logic;
  signal cond_br95_trueOut_valid : std_logic;
  signal cond_br95_trueOut_ready : std_logic;
  signal cond_br95_falseOut_valid : std_logic;
  signal cond_br95_falseOut_ready : std_logic;
  signal cond_br96_trueOut_valid : std_logic;
  signal cond_br96_trueOut_ready : std_logic;
  signal cond_br96_falseOut_valid : std_logic;
  signal cond_br96_falseOut_ready : std_logic;
  signal source13_outs_valid : std_logic;
  signal source13_outs_ready : std_logic;
  signal mux91_outs_valid : std_logic;
  signal mux91_outs_ready : std_logic;
  signal source14_outs_valid : std_logic;
  signal source14_outs_ready : std_logic;
  signal mux92_outs_valid : std_logic;
  signal mux92_outs_ready : std_logic;
  signal buffer50_outs_valid : std_logic;
  signal buffer50_outs_ready : std_logic;
  signal buffer51_outs_valid : std_logic;
  signal buffer51_outs_ready : std_logic;
  signal join3_outs_valid : std_logic;
  signal join3_outs_ready : std_logic;
  signal buffer52_outs_valid : std_logic;
  signal buffer52_outs_ready : std_logic;
  signal gate7_outs : std_logic_vector(31 downto 0);
  signal gate7_outs_valid : std_logic;
  signal gate7_outs_ready : std_logic;
  signal buffer148_outs : std_logic_vector(31 downto 0);
  signal buffer148_outs_valid : std_logic;
  signal buffer148_outs_ready : std_logic;
  signal trunci3_outs : std_logic_vector(6 downto 0);
  signal trunci3_outs_valid : std_logic;
  signal trunci3_outs_ready : std_logic;
  signal store0_addrOut : std_logic_vector(6 downto 0);
  signal store0_addrOut_valid : std_logic;
  signal store0_addrOut_ready : std_logic;
  signal store0_dataToMem : std_logic_vector(31 downto 0);
  signal store0_dataToMem_valid : std_logic;
  signal store0_dataToMem_ready : std_logic;
  signal store0_doneOut_valid : std_logic;
  signal store0_doneOut_ready : std_logic;
  signal addi4_result : std_logic_vector(8 downto 0);
  signal addi4_result_valid : std_logic;
  signal addi4_result_ready : std_logic;
  signal buffer54_outs : std_logic_vector(8 downto 0);
  signal buffer54_outs_valid : std_logic;
  signal buffer54_outs_ready : std_logic;
  signal fork50_outs_0 : std_logic_vector(8 downto 0);
  signal fork50_outs_0_valid : std_logic;
  signal fork50_outs_0_ready : std_logic;
  signal fork50_outs_1 : std_logic_vector(8 downto 0);
  signal fork50_outs_1_valid : std_logic;
  signal fork50_outs_1_ready : std_logic;
  signal trunci4_outs : std_logic_vector(7 downto 0);
  signal trunci4_outs_valid : std_logic;
  signal trunci4_outs_ready : std_logic;
  signal cmpi0_result : std_logic_vector(0 downto 0);
  signal cmpi0_result_valid : std_logic;
  signal cmpi0_result_ready : std_logic;
  signal fork51_outs_0 : std_logic_vector(0 downto 0);
  signal fork51_outs_0_valid : std_logic;
  signal fork51_outs_0_ready : std_logic;
  signal fork51_outs_1 : std_logic_vector(0 downto 0);
  signal fork51_outs_1_valid : std_logic;
  signal fork51_outs_1_ready : std_logic;
  signal fork51_outs_2 : std_logic_vector(0 downto 0);
  signal fork51_outs_2_valid : std_logic;
  signal fork51_outs_2_ready : std_logic;
  signal fork51_outs_3 : std_logic_vector(0 downto 0);
  signal fork51_outs_3_valid : std_logic;
  signal fork51_outs_3_ready : std_logic;
  signal fork51_outs_4 : std_logic_vector(0 downto 0);
  signal fork51_outs_4_valid : std_logic;
  signal fork51_outs_4_ready : std_logic;
  signal fork51_outs_5 : std_logic_vector(0 downto 0);
  signal fork51_outs_5_valid : std_logic;
  signal fork51_outs_5_ready : std_logic;
  signal fork51_outs_6 : std_logic_vector(0 downto 0);
  signal fork51_outs_6_valid : std_logic;
  signal fork51_outs_6_ready : std_logic;
  signal fork51_outs_7 : std_logic_vector(0 downto 0);
  signal fork51_outs_7_valid : std_logic;
  signal fork51_outs_7_ready : std_logic;
  signal fork51_outs_8 : std_logic_vector(0 downto 0);
  signal fork51_outs_8_valid : std_logic;
  signal fork51_outs_8_ready : std_logic;
  signal fork51_outs_9 : std_logic_vector(0 downto 0);
  signal fork51_outs_9_valid : std_logic;
  signal fork51_outs_9_ready : std_logic;
  signal fork51_outs_10 : std_logic_vector(0 downto 0);
  signal fork51_outs_10_valid : std_logic;
  signal fork51_outs_10_ready : std_logic;
  signal fork51_outs_11 : std_logic_vector(0 downto 0);
  signal fork51_outs_11_valid : std_logic;
  signal fork51_outs_11_ready : std_logic;
  signal fork51_outs_12 : std_logic_vector(0 downto 0);
  signal fork51_outs_12_valid : std_logic;
  signal fork51_outs_12_ready : std_logic;
  signal fork51_outs_13 : std_logic_vector(0 downto 0);
  signal fork51_outs_13_valid : std_logic;
  signal fork51_outs_13_ready : std_logic;
  signal fork51_outs_14 : std_logic_vector(0 downto 0);
  signal fork51_outs_14_valid : std_logic;
  signal fork51_outs_14_ready : std_logic;
  signal fork51_outs_15 : std_logic_vector(0 downto 0);
  signal fork51_outs_15_valid : std_logic;
  signal fork51_outs_15_ready : std_logic;
  signal fork51_outs_16 : std_logic_vector(0 downto 0);
  signal fork51_outs_16_valid : std_logic;
  signal fork51_outs_16_ready : std_logic;
  signal fork51_outs_17 : std_logic_vector(0 downto 0);
  signal fork51_outs_17_valid : std_logic;
  signal fork51_outs_17_ready : std_logic;
  signal fork51_outs_18 : std_logic_vector(0 downto 0);
  signal fork51_outs_18_valid : std_logic;
  signal fork51_outs_18_ready : std_logic;
  signal fork51_outs_19 : std_logic_vector(0 downto 0);
  signal fork51_outs_19_valid : std_logic;
  signal fork51_outs_19_ready : std_logic;
  signal fork51_outs_20 : std_logic_vector(0 downto 0);
  signal fork51_outs_20_valid : std_logic;
  signal fork51_outs_20_ready : std_logic;
  signal fork51_outs_21 : std_logic_vector(0 downto 0);
  signal fork51_outs_21_valid : std_logic;
  signal fork51_outs_21_ready : std_logic;
  signal fork51_outs_22 : std_logic_vector(0 downto 0);
  signal fork51_outs_22_valid : std_logic;
  signal fork51_outs_22_ready : std_logic;
  signal fork51_outs_23 : std_logic_vector(0 downto 0);
  signal fork51_outs_23_valid : std_logic;
  signal fork51_outs_23_ready : std_logic;
  signal fork51_outs_24 : std_logic_vector(0 downto 0);
  signal fork51_outs_24_valid : std_logic;
  signal fork51_outs_24_ready : std_logic;
  signal fork51_outs_25 : std_logic_vector(0 downto 0);
  signal fork51_outs_25_valid : std_logic;
  signal fork51_outs_25_ready : std_logic;
  signal fork51_outs_26 : std_logic_vector(0 downto 0);
  signal fork51_outs_26_valid : std_logic;
  signal fork51_outs_26_ready : std_logic;
  signal fork51_outs_27 : std_logic_vector(0 downto 0);
  signal fork51_outs_27_valid : std_logic;
  signal fork51_outs_27_ready : std_logic;
  signal fork51_outs_28 : std_logic_vector(0 downto 0);
  signal fork51_outs_28_valid : std_logic;
  signal fork51_outs_28_ready : std_logic;
  signal fork51_outs_29 : std_logic_vector(0 downto 0);
  signal fork51_outs_29_valid : std_logic;
  signal fork51_outs_29_ready : std_logic;
  signal fork51_outs_30 : std_logic_vector(0 downto 0);
  signal fork51_outs_30_valid : std_logic;
  signal fork51_outs_30_ready : std_logic;
  signal fork51_outs_31 : std_logic_vector(0 downto 0);
  signal fork51_outs_31_valid : std_logic;
  signal fork51_outs_31_ready : std_logic;
  signal fork51_outs_32 : std_logic_vector(0 downto 0);
  signal fork51_outs_32_valid : std_logic;
  signal fork51_outs_32_ready : std_logic;
  signal fork51_outs_33 : std_logic_vector(0 downto 0);
  signal fork51_outs_33_valid : std_logic;
  signal fork51_outs_33_ready : std_logic;
  signal cond_br3_trueOut : std_logic_vector(7 downto 0);
  signal cond_br3_trueOut_valid : std_logic;
  signal cond_br3_trueOut_ready : std_logic;
  signal cond_br3_falseOut : std_logic_vector(7 downto 0);
  signal cond_br3_falseOut_valid : std_logic;
  signal cond_br3_falseOut_ready : std_logic;
  signal buffer34_outs : std_logic_vector(2 downto 0);
  signal buffer34_outs_valid : std_logic;
  signal buffer34_outs_ready : std_logic;
  signal buffer35_outs : std_logic_vector(2 downto 0);
  signal buffer35_outs_valid : std_logic;
  signal buffer35_outs_ready : std_logic;
  signal cond_br4_trueOut : std_logic_vector(2 downto 0);
  signal cond_br4_trueOut_valid : std_logic;
  signal cond_br4_trueOut_ready : std_logic;
  signal cond_br4_falseOut : std_logic_vector(2 downto 0);
  signal cond_br4_falseOut_valid : std_logic;
  signal cond_br4_falseOut_ready : std_logic;
  signal cond_br5_trueOut_valid : std_logic;
  signal cond_br5_trueOut_ready : std_logic;
  signal cond_br5_falseOut_valid : std_logic;
  signal cond_br5_falseOut_ready : std_logic;
  signal cond_br6_trueOut : std_logic_vector(1 downto 0);
  signal cond_br6_trueOut_valid : std_logic;
  signal cond_br6_trueOut_ready : std_logic;
  signal cond_br6_falseOut : std_logic_vector(1 downto 0);
  signal cond_br6_falseOut_valid : std_logic;
  signal cond_br6_falseOut_ready : std_logic;
  signal extsi19_outs : std_logic_vector(7 downto 0);
  signal extsi19_outs_valid : std_logic;
  signal extsi19_outs_ready : std_logic;
  signal cond_br234_trueOut : std_logic_vector(8 downto 0);
  signal cond_br234_trueOut_valid : std_logic;
  signal cond_br234_trueOut_ready : std_logic;
  signal cond_br234_falseOut : std_logic_vector(8 downto 0);
  signal cond_br234_falseOut_valid : std_logic;
  signal cond_br234_falseOut_ready : std_logic;
  signal cond_br235_trueOut : std_logic_vector(31 downto 0);
  signal cond_br235_trueOut_valid : std_logic;
  signal cond_br235_trueOut_ready : std_logic;
  signal cond_br235_falseOut : std_logic_vector(31 downto 0);
  signal cond_br235_falseOut_valid : std_logic;
  signal cond_br235_falseOut_ready : std_logic;
  signal cond_br236_trueOut_valid : std_logic;
  signal cond_br236_trueOut_ready : std_logic;
  signal cond_br236_falseOut_valid : std_logic;
  signal cond_br236_falseOut_ready : std_logic;
  signal buffer160_outs : std_logic_vector(0 downto 0);
  signal buffer160_outs_valid : std_logic;
  signal buffer160_outs_ready : std_logic;
  signal cond_br237_trueOut_valid : std_logic;
  signal cond_br237_trueOut_ready : std_logic;
  signal cond_br237_falseOut_valid : std_logic;
  signal cond_br237_falseOut_ready : std_logic;
  signal cond_br238_trueOut_valid : std_logic;
  signal cond_br238_trueOut_ready : std_logic;
  signal cond_br238_falseOut_valid : std_logic;
  signal cond_br238_falseOut_ready : std_logic;
  signal cond_br239_trueOut : std_logic_vector(31 downto 0);
  signal cond_br239_trueOut_valid : std_logic;
  signal cond_br239_trueOut_ready : std_logic;
  signal cond_br239_falseOut : std_logic_vector(31 downto 0);
  signal cond_br239_falseOut_valid : std_logic;
  signal cond_br239_falseOut_ready : std_logic;
  signal cond_br240_trueOut_valid : std_logic;
  signal cond_br240_trueOut_ready : std_logic;
  signal cond_br240_falseOut_valid : std_logic;
  signal cond_br240_falseOut_ready : std_logic;
  signal cond_br241_trueOut_valid : std_logic;
  signal cond_br241_trueOut_ready : std_logic;
  signal cond_br241_falseOut_valid : std_logic;
  signal cond_br241_falseOut_ready : std_logic;
  signal cond_br242_trueOut : std_logic_vector(7 downto 0);
  signal cond_br242_trueOut_valid : std_logic;
  signal cond_br242_trueOut_ready : std_logic;
  signal cond_br242_falseOut : std_logic_vector(7 downto 0);
  signal cond_br242_falseOut_valid : std_logic;
  signal cond_br242_falseOut_ready : std_logic;
  signal cond_br243_trueOut_valid : std_logic;
  signal cond_br243_trueOut_ready : std_logic;
  signal cond_br243_falseOut_valid : std_logic;
  signal cond_br243_falseOut_ready : std_logic;
  signal cond_br244_trueOut : std_logic_vector(31 downto 0);
  signal cond_br244_trueOut_valid : std_logic;
  signal cond_br244_trueOut_ready : std_logic;
  signal cond_br244_falseOut : std_logic_vector(31 downto 0);
  signal cond_br244_falseOut_valid : std_logic;
  signal cond_br244_falseOut_ready : std_logic;
  signal cond_br245_trueOut_valid : std_logic;
  signal cond_br245_trueOut_ready : std_logic;
  signal cond_br245_falseOut_valid : std_logic;
  signal cond_br245_falseOut_ready : std_logic;
  signal cond_br246_trueOut : std_logic_vector(7 downto 0);
  signal cond_br246_trueOut_valid : std_logic;
  signal cond_br246_trueOut_ready : std_logic;
  signal cond_br246_falseOut : std_logic_vector(7 downto 0);
  signal cond_br246_falseOut_valid : std_logic;
  signal cond_br246_falseOut_ready : std_logic;
  signal cond_br247_trueOut_valid : std_logic;
  signal cond_br247_trueOut_ready : std_logic;
  signal cond_br247_falseOut_valid : std_logic;
  signal cond_br247_falseOut_ready : std_logic;
  signal buffer174_outs : std_logic_vector(0 downto 0);
  signal buffer174_outs_valid : std_logic;
  signal buffer174_outs_ready : std_logic;
  signal cond_br248_trueOut_valid : std_logic;
  signal cond_br248_trueOut_ready : std_logic;
  signal cond_br248_falseOut_valid : std_logic;
  signal cond_br248_falseOut_ready : std_logic;
  signal buffer175_outs : std_logic_vector(0 downto 0);
  signal buffer175_outs_valid : std_logic;
  signal buffer175_outs_ready : std_logic;
  signal cond_br249_trueOut : std_logic_vector(31 downto 0);
  signal cond_br249_trueOut_valid : std_logic;
  signal cond_br249_trueOut_ready : std_logic;
  signal cond_br249_falseOut : std_logic_vector(31 downto 0);
  signal cond_br249_falseOut_valid : std_logic;
  signal cond_br249_falseOut_ready : std_logic;
  signal cond_br250_trueOut_valid : std_logic;
  signal cond_br250_trueOut_ready : std_logic;
  signal cond_br250_falseOut_valid : std_logic;
  signal cond_br250_falseOut_ready : std_logic;
  signal buffer177_outs : std_logic_vector(0 downto 0);
  signal buffer177_outs_valid : std_logic;
  signal buffer177_outs_ready : std_logic;
  signal cond_br251_trueOut : std_logic_vector(31 downto 0);
  signal cond_br251_trueOut_valid : std_logic;
  signal cond_br251_trueOut_ready : std_logic;
  signal cond_br251_falseOut : std_logic_vector(31 downto 0);
  signal cond_br251_falseOut_valid : std_logic;
  signal cond_br251_falseOut_ready : std_logic;
  signal buffer179_outs : std_logic_vector(31 downto 0);
  signal buffer179_outs_valid : std_logic;
  signal buffer179_outs_ready : std_logic;
  signal cond_br252_trueOut : std_logic_vector(7 downto 0);
  signal cond_br252_trueOut_valid : std_logic;
  signal cond_br252_trueOut_ready : std_logic;
  signal cond_br252_falseOut : std_logic_vector(7 downto 0);
  signal cond_br252_falseOut_valid : std_logic;
  signal cond_br252_falseOut_ready : std_logic;
  signal buffer180_outs : std_logic_vector(0 downto 0);
  signal buffer180_outs_valid : std_logic;
  signal buffer180_outs_ready : std_logic;
  signal cond_br253_trueOut_valid : std_logic;
  signal cond_br253_trueOut_ready : std_logic;
  signal cond_br253_falseOut_valid : std_logic;
  signal cond_br253_falseOut_ready : std_logic;
  signal cond_br254_trueOut : std_logic_vector(31 downto 0);
  signal cond_br254_trueOut_valid : std_logic;
  signal cond_br254_trueOut_ready : std_logic;
  signal cond_br254_falseOut : std_logic_vector(31 downto 0);
  signal cond_br254_falseOut_valid : std_logic;
  signal cond_br254_falseOut_ready : std_logic;
  signal buffer184_outs : std_logic_vector(31 downto 0);
  signal buffer184_outs_valid : std_logic;
  signal buffer184_outs_ready : std_logic;
  signal cond_br255_trueOut_valid : std_logic;
  signal cond_br255_trueOut_ready : std_logic;
  signal cond_br255_falseOut_valid : std_logic;
  signal cond_br255_falseOut_ready : std_logic;
  signal buffer185_outs : std_logic_vector(0 downto 0);
  signal buffer185_outs_valid : std_logic;
  signal buffer185_outs_ready : std_logic;
  signal cond_br256_trueOut : std_logic_vector(31 downto 0);
  signal cond_br256_trueOut_valid : std_logic;
  signal cond_br256_trueOut_ready : std_logic;
  signal cond_br256_falseOut : std_logic_vector(31 downto 0);
  signal cond_br256_falseOut_valid : std_logic;
  signal cond_br256_falseOut_ready : std_logic;
  signal buffer186_outs : std_logic_vector(0 downto 0);
  signal buffer186_outs_valid : std_logic;
  signal buffer186_outs_ready : std_logic;
  signal buffer187_outs : std_logic_vector(31 downto 0);
  signal buffer187_outs_valid : std_logic;
  signal buffer187_outs_ready : std_logic;
  signal cond_br257_trueOut_valid : std_logic;
  signal cond_br257_trueOut_ready : std_logic;
  signal cond_br257_falseOut_valid : std_logic;
  signal cond_br257_falseOut_ready : std_logic;
  signal buffer188_outs : std_logic_vector(0 downto 0);
  signal buffer188_outs_valid : std_logic;
  signal buffer188_outs_ready : std_logic;
  signal cond_br258_trueOut : std_logic_vector(7 downto 0);
  signal cond_br258_trueOut_valid : std_logic;
  signal cond_br258_trueOut_ready : std_logic;
  signal cond_br258_falseOut : std_logic_vector(7 downto 0);
  signal cond_br258_falseOut_valid : std_logic;
  signal cond_br258_falseOut_ready : std_logic;
  signal init92_outs : std_logic_vector(0 downto 0);
  signal init92_outs_valid : std_logic;
  signal init92_outs_ready : std_logic;
  signal fork52_outs_0 : std_logic_vector(0 downto 0);
  signal fork52_outs_0_valid : std_logic;
  signal fork52_outs_0_ready : std_logic;
  signal fork52_outs_1 : std_logic_vector(0 downto 0);
  signal fork52_outs_1_valid : std_logic;
  signal fork52_outs_1_ready : std_logic;
  signal fork52_outs_2 : std_logic_vector(0 downto 0);
  signal fork52_outs_2_valid : std_logic;
  signal fork52_outs_2_ready : std_logic;
  signal fork52_outs_3 : std_logic_vector(0 downto 0);
  signal fork52_outs_3_valid : std_logic;
  signal fork52_outs_3_ready : std_logic;
  signal fork52_outs_4 : std_logic_vector(0 downto 0);
  signal fork52_outs_4_valid : std_logic;
  signal fork52_outs_4_ready : std_logic;
  signal fork52_outs_5 : std_logic_vector(0 downto 0);
  signal fork52_outs_5_valid : std_logic;
  signal fork52_outs_5_ready : std_logic;
  signal fork52_outs_6 : std_logic_vector(0 downto 0);
  signal fork52_outs_6_valid : std_logic;
  signal fork52_outs_6_ready : std_logic;
  signal fork52_outs_7 : std_logic_vector(0 downto 0);
  signal fork52_outs_7_valid : std_logic;
  signal fork52_outs_7_ready : std_logic;
  signal fork52_outs_8 : std_logic_vector(0 downto 0);
  signal fork52_outs_8_valid : std_logic;
  signal fork52_outs_8_ready : std_logic;
  signal fork52_outs_9 : std_logic_vector(0 downto 0);
  signal fork52_outs_9_valid : std_logic;
  signal fork52_outs_9_ready : std_logic;
  signal fork52_outs_10 : std_logic_vector(0 downto 0);
  signal fork52_outs_10_valid : std_logic;
  signal fork52_outs_10_ready : std_logic;
  signal fork52_outs_11 : std_logic_vector(0 downto 0);
  signal fork52_outs_11_valid : std_logic;
  signal fork52_outs_11_ready : std_logic;
  signal fork52_outs_12 : std_logic_vector(0 downto 0);
  signal fork52_outs_12_valid : std_logic;
  signal fork52_outs_12_ready : std_logic;
  signal fork52_outs_13 : std_logic_vector(0 downto 0);
  signal fork52_outs_13_valid : std_logic;
  signal fork52_outs_13_ready : std_logic;
  signal fork52_outs_14 : std_logic_vector(0 downto 0);
  signal fork52_outs_14_valid : std_logic;
  signal fork52_outs_14_ready : std_logic;
  signal fork52_outs_15 : std_logic_vector(0 downto 0);
  signal fork52_outs_15_valid : std_logic;
  signal fork52_outs_15_ready : std_logic;
  signal fork52_outs_16 : std_logic_vector(0 downto 0);
  signal fork52_outs_16_valid : std_logic;
  signal fork52_outs_16_ready : std_logic;
  signal fork52_outs_17 : std_logic_vector(0 downto 0);
  signal fork52_outs_17_valid : std_logic;
  signal fork52_outs_17_ready : std_logic;
  signal fork52_outs_18 : std_logic_vector(0 downto 0);
  signal fork52_outs_18_valid : std_logic;
  signal fork52_outs_18_ready : std_logic;
  signal fork52_outs_19 : std_logic_vector(0 downto 0);
  signal fork52_outs_19_valid : std_logic;
  signal fork52_outs_19_ready : std_logic;
  signal mux93_outs : std_logic_vector(7 downto 0);
  signal mux93_outs_valid : std_logic;
  signal mux93_outs_ready : std_logic;
  signal buffer55_outs : std_logic_vector(7 downto 0);
  signal buffer55_outs_valid : std_logic;
  signal buffer55_outs_ready : std_logic;
  signal buffer56_outs : std_logic_vector(7 downto 0);
  signal buffer56_outs_valid : std_logic;
  signal buffer56_outs_ready : std_logic;
  signal fork53_outs_0 : std_logic_vector(7 downto 0);
  signal fork53_outs_0_valid : std_logic;
  signal fork53_outs_0_ready : std_logic;
  signal fork53_outs_1 : std_logic_vector(7 downto 0);
  signal fork53_outs_1_valid : std_logic;
  signal fork53_outs_1_ready : std_logic;
  signal extsi36_outs : std_logic_vector(31 downto 0);
  signal extsi36_outs_valid : std_logic;
  signal extsi36_outs_ready : std_logic;
  signal buffer193_outs : std_logic_vector(7 downto 0);
  signal buffer193_outs_valid : std_logic;
  signal buffer193_outs_ready : std_logic;
  signal mux94_outs_valid : std_logic;
  signal mux94_outs_ready : std_logic;
  signal buffer194_outs : std_logic_vector(0 downto 0);
  signal buffer194_outs_valid : std_logic;
  signal buffer194_outs_ready : std_logic;
  signal buffer58_outs_valid : std_logic;
  signal buffer58_outs_ready : std_logic;
  signal buffer59_outs_valid : std_logic;
  signal buffer59_outs_ready : std_logic;
  signal fork54_outs_0_valid : std_logic;
  signal fork54_outs_0_ready : std_logic;
  signal fork54_outs_1_valid : std_logic;
  signal fork54_outs_1_ready : std_logic;
  signal mux95_outs : std_logic_vector(31 downto 0);
  signal mux95_outs_valid : std_logic;
  signal mux95_outs_ready : std_logic;
  signal buffer195_outs : std_logic_vector(0 downto 0);
  signal buffer195_outs_valid : std_logic;
  signal buffer195_outs_ready : std_logic;
  signal buffer60_outs : std_logic_vector(31 downto 0);
  signal buffer60_outs_valid : std_logic;
  signal buffer60_outs_ready : std_logic;
  signal buffer61_outs : std_logic_vector(31 downto 0);
  signal buffer61_outs_valid : std_logic;
  signal buffer61_outs_ready : std_logic;
  signal fork55_outs_0 : std_logic_vector(31 downto 0);
  signal fork55_outs_0_valid : std_logic;
  signal fork55_outs_0_ready : std_logic;
  signal fork55_outs_1 : std_logic_vector(31 downto 0);
  signal fork55_outs_1_valid : std_logic;
  signal fork55_outs_1_ready : std_logic;
  signal mux96_outs_valid : std_logic;
  signal mux96_outs_ready : std_logic;
  signal buffer196_outs : std_logic_vector(0 downto 0);
  signal buffer196_outs_valid : std_logic;
  signal buffer196_outs_ready : std_logic;
  signal buffer62_outs_valid : std_logic;
  signal buffer62_outs_ready : std_logic;
  signal buffer63_outs_valid : std_logic;
  signal buffer63_outs_ready : std_logic;
  signal fork56_outs_0_valid : std_logic;
  signal fork56_outs_0_ready : std_logic;
  signal fork56_outs_1_valid : std_logic;
  signal fork56_outs_1_ready : std_logic;
  signal mux97_outs : std_logic_vector(8 downto 0);
  signal mux97_outs_valid : std_logic;
  signal mux97_outs_ready : std_logic;
  signal buffer197_outs : std_logic_vector(0 downto 0);
  signal buffer197_outs_valid : std_logic;
  signal buffer197_outs_ready : std_logic;
  signal buffer64_outs : std_logic_vector(8 downto 0);
  signal buffer64_outs_valid : std_logic;
  signal buffer64_outs_ready : std_logic;
  signal buffer65_outs : std_logic_vector(8 downto 0);
  signal buffer65_outs_valid : std_logic;
  signal buffer65_outs_ready : std_logic;
  signal fork57_outs_0 : std_logic_vector(8 downto 0);
  signal fork57_outs_0_valid : std_logic;
  signal fork57_outs_0_ready : std_logic;
  signal fork57_outs_1 : std_logic_vector(8 downto 0);
  signal fork57_outs_1_valid : std_logic;
  signal fork57_outs_1_ready : std_logic;
  signal extsi37_outs : std_logic_vector(31 downto 0);
  signal extsi37_outs_valid : std_logic;
  signal extsi37_outs_ready : std_logic;
  signal buffer198_outs : std_logic_vector(8 downto 0);
  signal buffer198_outs_valid : std_logic;
  signal buffer198_outs_ready : std_logic;
  signal mux98_outs : std_logic_vector(7 downto 0);
  signal mux98_outs_valid : std_logic;
  signal mux98_outs_ready : std_logic;
  signal buffer199_outs : std_logic_vector(0 downto 0);
  signal buffer199_outs_valid : std_logic;
  signal buffer199_outs_ready : std_logic;
  signal buffer67_outs : std_logic_vector(7 downto 0);
  signal buffer67_outs_valid : std_logic;
  signal buffer67_outs_ready : std_logic;
  signal buffer69_outs : std_logic_vector(7 downto 0);
  signal buffer69_outs_valid : std_logic;
  signal buffer69_outs_ready : std_logic;
  signal fork58_outs_0 : std_logic_vector(7 downto 0);
  signal fork58_outs_0_valid : std_logic;
  signal fork58_outs_0_ready : std_logic;
  signal fork58_outs_1 : std_logic_vector(7 downto 0);
  signal fork58_outs_1_valid : std_logic;
  signal fork58_outs_1_ready : std_logic;
  signal extsi38_outs : std_logic_vector(31 downto 0);
  signal extsi38_outs_valid : std_logic;
  signal extsi38_outs_ready : std_logic;
  signal buffer200_outs : std_logic_vector(7 downto 0);
  signal buffer200_outs_valid : std_logic;
  signal buffer200_outs_ready : std_logic;
  signal mux99_outs : std_logic_vector(31 downto 0);
  signal mux99_outs_valid : std_logic;
  signal mux99_outs_ready : std_logic;
  signal buffer201_outs : std_logic_vector(0 downto 0);
  signal buffer201_outs_valid : std_logic;
  signal buffer201_outs_ready : std_logic;
  signal buffer70_outs : std_logic_vector(31 downto 0);
  signal buffer70_outs_valid : std_logic;
  signal buffer70_outs_ready : std_logic;
  signal buffer71_outs : std_logic_vector(31 downto 0);
  signal buffer71_outs_valid : std_logic;
  signal buffer71_outs_ready : std_logic;
  signal fork59_outs_0 : std_logic_vector(31 downto 0);
  signal fork59_outs_0_valid : std_logic;
  signal fork59_outs_0_ready : std_logic;
  signal fork59_outs_1 : std_logic_vector(31 downto 0);
  signal fork59_outs_1_valid : std_logic;
  signal fork59_outs_1_ready : std_logic;
  signal mux100_outs_valid : std_logic;
  signal mux100_outs_ready : std_logic;
  signal buffer202_outs : std_logic_vector(0 downto 0);
  signal buffer202_outs_valid : std_logic;
  signal buffer202_outs_ready : std_logic;
  signal buffer72_outs_valid : std_logic;
  signal buffer72_outs_ready : std_logic;
  signal buffer73_outs_valid : std_logic;
  signal buffer73_outs_ready : std_logic;
  signal fork60_outs_0_valid : std_logic;
  signal fork60_outs_0_ready : std_logic;
  signal fork60_outs_1_valid : std_logic;
  signal fork60_outs_1_ready : std_logic;
  signal mux101_outs_valid : std_logic;
  signal mux101_outs_ready : std_logic;
  signal buffer203_outs : std_logic_vector(0 downto 0);
  signal buffer203_outs_valid : std_logic;
  signal buffer203_outs_ready : std_logic;
  signal buffer74_outs_valid : std_logic;
  signal buffer74_outs_ready : std_logic;
  signal buffer75_outs_valid : std_logic;
  signal buffer75_outs_ready : std_logic;
  signal fork61_outs_0_valid : std_logic;
  signal fork61_outs_0_ready : std_logic;
  signal fork61_outs_1_valid : std_logic;
  signal fork61_outs_1_ready : std_logic;
  signal mux102_outs_valid : std_logic;
  signal mux102_outs_ready : std_logic;
  signal buffer204_outs : std_logic_vector(0 downto 0);
  signal buffer204_outs_valid : std_logic;
  signal buffer204_outs_ready : std_logic;
  signal buffer76_outs_valid : std_logic;
  signal buffer76_outs_ready : std_logic;
  signal buffer77_outs_valid : std_logic;
  signal buffer77_outs_ready : std_logic;
  signal fork62_outs_0_valid : std_logic;
  signal fork62_outs_0_ready : std_logic;
  signal fork62_outs_1_valid : std_logic;
  signal fork62_outs_1_ready : std_logic;
  signal mux103_outs : std_logic_vector(31 downto 0);
  signal mux103_outs_valid : std_logic;
  signal mux103_outs_ready : std_logic;
  signal buffer205_outs : std_logic_vector(0 downto 0);
  signal buffer205_outs_valid : std_logic;
  signal buffer205_outs_ready : std_logic;
  signal buffer78_outs : std_logic_vector(31 downto 0);
  signal buffer78_outs_valid : std_logic;
  signal buffer78_outs_ready : std_logic;
  signal buffer79_outs : std_logic_vector(31 downto 0);
  signal buffer79_outs_valid : std_logic;
  signal buffer79_outs_ready : std_logic;
  signal fork63_outs_0 : std_logic_vector(31 downto 0);
  signal fork63_outs_0_valid : std_logic;
  signal fork63_outs_0_ready : std_logic;
  signal fork63_outs_1 : std_logic_vector(31 downto 0);
  signal fork63_outs_1_valid : std_logic;
  signal fork63_outs_1_ready : std_logic;
  signal mux104_outs_valid : std_logic;
  signal mux104_outs_ready : std_logic;
  signal buffer206_outs : std_logic_vector(0 downto 0);
  signal buffer206_outs_valid : std_logic;
  signal buffer206_outs_ready : std_logic;
  signal buffer80_outs_valid : std_logic;
  signal buffer80_outs_ready : std_logic;
  signal buffer81_outs_valid : std_logic;
  signal buffer81_outs_ready : std_logic;
  signal fork64_outs_0_valid : std_logic;
  signal fork64_outs_0_ready : std_logic;
  signal fork64_outs_1_valid : std_logic;
  signal fork64_outs_1_ready : std_logic;
  signal mux105_outs_valid : std_logic;
  signal mux105_outs_ready : std_logic;
  signal buffer207_outs : std_logic_vector(0 downto 0);
  signal buffer207_outs_valid : std_logic;
  signal buffer207_outs_ready : std_logic;
  signal buffer82_outs_valid : std_logic;
  signal buffer82_outs_ready : std_logic;
  signal buffer83_outs_valid : std_logic;
  signal buffer83_outs_ready : std_logic;
  signal fork65_outs_0_valid : std_logic;
  signal fork65_outs_0_ready : std_logic;
  signal fork65_outs_1_valid : std_logic;
  signal fork65_outs_1_ready : std_logic;
  signal mux106_outs_valid : std_logic;
  signal mux106_outs_ready : std_logic;
  signal buffer84_outs_valid : std_logic;
  signal buffer84_outs_ready : std_logic;
  signal buffer85_outs_valid : std_logic;
  signal buffer85_outs_ready : std_logic;
  signal fork66_outs_0_valid : std_logic;
  signal fork66_outs_0_ready : std_logic;
  signal fork66_outs_1_valid : std_logic;
  signal fork66_outs_1_ready : std_logic;
  signal mux107_outs_valid : std_logic;
  signal mux107_outs_ready : std_logic;
  signal buffer209_outs : std_logic_vector(0 downto 0);
  signal buffer209_outs_valid : std_logic;
  signal buffer209_outs_ready : std_logic;
  signal buffer86_outs_valid : std_logic;
  signal buffer86_outs_ready : std_logic;
  signal buffer87_outs_valid : std_logic;
  signal buffer87_outs_ready : std_logic;
  signal fork67_outs_0_valid : std_logic;
  signal fork67_outs_0_ready : std_logic;
  signal fork67_outs_1_valid : std_logic;
  signal fork67_outs_1_ready : std_logic;
  signal mux108_outs_valid : std_logic;
  signal mux108_outs_ready : std_logic;
  signal buffer210_outs : std_logic_vector(0 downto 0);
  signal buffer210_outs_valid : std_logic;
  signal buffer210_outs_ready : std_logic;
  signal buffer88_outs_valid : std_logic;
  signal buffer88_outs_ready : std_logic;
  signal buffer89_outs_valid : std_logic;
  signal buffer89_outs_ready : std_logic;
  signal fork68_outs_0_valid : std_logic;
  signal fork68_outs_0_ready : std_logic;
  signal fork68_outs_1_valid : std_logic;
  signal fork68_outs_1_ready : std_logic;
  signal mux109_outs : std_logic_vector(31 downto 0);
  signal mux109_outs_valid : std_logic;
  signal mux109_outs_ready : std_logic;
  signal buffer211_outs : std_logic_vector(0 downto 0);
  signal buffer211_outs_valid : std_logic;
  signal buffer211_outs_ready : std_logic;
  signal buffer90_outs : std_logic_vector(31 downto 0);
  signal buffer90_outs_valid : std_logic;
  signal buffer90_outs_ready : std_logic;
  signal buffer91_outs : std_logic_vector(31 downto 0);
  signal buffer91_outs_valid : std_logic;
  signal buffer91_outs_ready : std_logic;
  signal fork69_outs_0 : std_logic_vector(31 downto 0);
  signal fork69_outs_0_valid : std_logic;
  signal fork69_outs_0_ready : std_logic;
  signal fork69_outs_1 : std_logic_vector(31 downto 0);
  signal fork69_outs_1_valid : std_logic;
  signal fork69_outs_1_ready : std_logic;
  signal mux110_outs : std_logic_vector(31 downto 0);
  signal mux110_outs_valid : std_logic;
  signal mux110_outs_ready : std_logic;
  signal buffer212_outs : std_logic_vector(0 downto 0);
  signal buffer212_outs_valid : std_logic;
  signal buffer212_outs_ready : std_logic;
  signal buffer92_outs : std_logic_vector(31 downto 0);
  signal buffer92_outs_valid : std_logic;
  signal buffer92_outs_ready : std_logic;
  signal buffer93_outs : std_logic_vector(31 downto 0);
  signal buffer93_outs_valid : std_logic;
  signal buffer93_outs_ready : std_logic;
  signal fork70_outs_0 : std_logic_vector(31 downto 0);
  signal fork70_outs_0_valid : std_logic;
  signal fork70_outs_0_ready : std_logic;
  signal fork70_outs_1 : std_logic_vector(31 downto 0);
  signal fork70_outs_1_valid : std_logic;
  signal fork70_outs_1_ready : std_logic;
  signal mux111_outs_valid : std_logic;
  signal mux111_outs_ready : std_logic;
  signal buffer213_outs : std_logic_vector(0 downto 0);
  signal buffer213_outs_valid : std_logic;
  signal buffer213_outs_ready : std_logic;
  signal buffer94_outs_valid : std_logic;
  signal buffer94_outs_ready : std_logic;
  signal buffer95_outs_valid : std_logic;
  signal buffer95_outs_ready : std_logic;
  signal fork71_outs_0_valid : std_logic;
  signal fork71_outs_0_ready : std_logic;
  signal fork71_outs_1_valid : std_logic;
  signal fork71_outs_1_ready : std_logic;
  signal mux112_outs_valid : std_logic;
  signal mux112_outs_ready : std_logic;
  signal buffer214_outs : std_logic_vector(0 downto 0);
  signal buffer214_outs_valid : std_logic;
  signal buffer214_outs_ready : std_logic;
  signal buffer96_outs_valid : std_logic;
  signal buffer96_outs_ready : std_logic;
  signal buffer97_outs_valid : std_logic;
  signal buffer97_outs_ready : std_logic;
  signal fork72_outs_0_valid : std_logic;
  signal fork72_outs_0_ready : std_logic;
  signal fork72_outs_1_valid : std_logic;
  signal fork72_outs_1_ready : std_logic;
  signal unbundle7_outs_0_valid : std_logic;
  signal unbundle7_outs_0_ready : std_logic;
  signal unbundle7_outs_1 : std_logic_vector(31 downto 0);
  signal mux3_outs : std_logic_vector(7 downto 0);
  signal mux3_outs_valid : std_logic;
  signal mux3_outs_ready : std_logic;
  signal buffer98_outs : std_logic_vector(7 downto 0);
  signal buffer98_outs_valid : std_logic;
  signal buffer98_outs_ready : std_logic;
  signal buffer99_outs : std_logic_vector(7 downto 0);
  signal buffer99_outs_valid : std_logic;
  signal buffer99_outs_ready : std_logic;
  signal fork73_outs_0 : std_logic_vector(7 downto 0);
  signal fork73_outs_0_valid : std_logic;
  signal fork73_outs_0_ready : std_logic;
  signal fork73_outs_1 : std_logic_vector(7 downto 0);
  signal fork73_outs_1_valid : std_logic;
  signal fork73_outs_1_ready : std_logic;
  signal fork73_outs_2 : std_logic_vector(7 downto 0);
  signal fork73_outs_2_valid : std_logic;
  signal fork73_outs_2_ready : std_logic;
  signal fork73_outs_3 : std_logic_vector(7 downto 0);
  signal fork73_outs_3_valid : std_logic;
  signal fork73_outs_3_ready : std_logic;
  signal extsi39_outs : std_logic_vector(8 downto 0);
  signal extsi39_outs_valid : std_logic;
  signal extsi39_outs_ready : std_logic;
  signal extsi40_outs : std_logic_vector(31 downto 0);
  signal extsi40_outs_valid : std_logic;
  signal extsi40_outs_ready : std_logic;
  signal buffer218_outs : std_logic_vector(7 downto 0);
  signal buffer218_outs_valid : std_logic;
  signal buffer218_outs_ready : std_logic;
  signal fork74_outs_0 : std_logic_vector(31 downto 0);
  signal fork74_outs_0_valid : std_logic;
  signal fork74_outs_0_ready : std_logic;
  signal fork74_outs_1 : std_logic_vector(31 downto 0);
  signal fork74_outs_1_valid : std_logic;
  signal fork74_outs_1_ready : std_logic;
  signal fork74_outs_2 : std_logic_vector(31 downto 0);
  signal fork74_outs_2_valid : std_logic;
  signal fork74_outs_2_ready : std_logic;
  signal fork74_outs_3 : std_logic_vector(31 downto 0);
  signal fork74_outs_3_valid : std_logic;
  signal fork74_outs_3_ready : std_logic;
  signal fork74_outs_4 : std_logic_vector(31 downto 0);
  signal fork74_outs_4_valid : std_logic;
  signal fork74_outs_4_ready : std_logic;
  signal fork74_outs_5 : std_logic_vector(31 downto 0);
  signal fork74_outs_5_valid : std_logic;
  signal fork74_outs_5_ready : std_logic;
  signal mux4_outs : std_logic_vector(2 downto 0);
  signal mux4_outs_valid : std_logic;
  signal mux4_outs_ready : std_logic;
  signal control_merge2_outs_valid : std_logic;
  signal control_merge2_outs_ready : std_logic;
  signal control_merge2_index : std_logic_vector(0 downto 0);
  signal control_merge2_index_valid : std_logic;
  signal control_merge2_index_ready : std_logic;
  signal fork75_outs_0 : std_logic_vector(0 downto 0);
  signal fork75_outs_0_valid : std_logic;
  signal fork75_outs_0_ready : std_logic;
  signal fork75_outs_1 : std_logic_vector(0 downto 0);
  signal fork75_outs_1_valid : std_logic;
  signal fork75_outs_1_ready : std_logic;
  signal fork76_outs_0_valid : std_logic;
  signal fork76_outs_0_ready : std_logic;
  signal fork76_outs_1_valid : std_logic;
  signal fork76_outs_1_ready : std_logic;
  signal constant20_outs : std_logic_vector(1 downto 0);
  signal constant20_outs_valid : std_logic;
  signal constant20_outs_ready : std_logic;
  signal extsi14_outs : std_logic_vector(31 downto 0);
  signal extsi14_outs_valid : std_logic;
  signal extsi14_outs_ready : std_logic;
  signal source3_outs_valid : std_logic;
  signal source3_outs_ready : std_logic;
  signal constant25_outs : std_logic_vector(7 downto 0);
  signal constant25_outs_valid : std_logic;
  signal constant25_outs_ready : std_logic;
  signal extsi41_outs : std_logic_vector(8 downto 0);
  signal extsi41_outs_valid : std_logic;
  signal extsi41_outs_ready : std_logic;
  signal source4_outs_valid : std_logic;
  signal source4_outs_ready : std_logic;
  signal constant28_outs : std_logic_vector(1 downto 0);
  signal constant28_outs_valid : std_logic;
  signal constant28_outs_ready : std_logic;
  signal extsi42_outs : std_logic_vector(8 downto 0);
  signal extsi42_outs_valid : std_logic;
  signal extsi42_outs_ready : std_logic;
  signal gate8_outs : std_logic_vector(31 downto 0);
  signal gate8_outs_valid : std_logic;
  signal gate8_outs_ready : std_logic;
  signal buffer220_outs : std_logic_vector(31 downto 0);
  signal buffer220_outs_valid : std_logic;
  signal buffer220_outs_ready : std_logic;
  signal fork77_outs_0 : std_logic_vector(31 downto 0);
  signal fork77_outs_0_valid : std_logic;
  signal fork77_outs_0_ready : std_logic;
  signal fork77_outs_1 : std_logic_vector(31 downto 0);
  signal fork77_outs_1_valid : std_logic;
  signal fork77_outs_1_ready : std_logic;
  signal cmpi11_result : std_logic_vector(0 downto 0);
  signal cmpi11_result_valid : std_logic;
  signal cmpi11_result_ready : std_logic;
  signal fork78_outs_0 : std_logic_vector(0 downto 0);
  signal fork78_outs_0_valid : std_logic;
  signal fork78_outs_0_ready : std_logic;
  signal fork78_outs_1 : std_logic_vector(0 downto 0);
  signal fork78_outs_1_valid : std_logic;
  signal fork78_outs_1_ready : std_logic;
  signal cmpi12_result : std_logic_vector(0 downto 0);
  signal cmpi12_result_valid : std_logic;
  signal cmpi12_result_ready : std_logic;
  signal buffer223_outs : std_logic_vector(31 downto 0);
  signal buffer223_outs_valid : std_logic;
  signal buffer223_outs_ready : std_logic;
  signal fork79_outs_0 : std_logic_vector(0 downto 0);
  signal fork79_outs_0_valid : std_logic;
  signal fork79_outs_0_ready : std_logic;
  signal fork79_outs_1 : std_logic_vector(0 downto 0);
  signal fork79_outs_1_valid : std_logic;
  signal fork79_outs_1_ready : std_logic;
  signal buffer8_outs : std_logic_vector(7 downto 0);
  signal buffer8_outs_valid : std_logic;
  signal buffer8_outs_ready : std_logic;
  signal fork80_outs_0 : std_logic_vector(7 downto 0);
  signal fork80_outs_0_valid : std_logic;
  signal fork80_outs_0_ready : std_logic;
  signal fork80_outs_1 : std_logic_vector(7 downto 0);
  signal fork80_outs_1_valid : std_logic;
  signal fork80_outs_1_ready : std_logic;
  signal extsi43_outs : std_logic_vector(31 downto 0);
  signal extsi43_outs_valid : std_logic;
  signal extsi43_outs_ready : std_logic;
  signal buffer225_outs : std_logic_vector(7 downto 0);
  signal buffer225_outs_valid : std_logic;
  signal buffer225_outs_ready : std_logic;
  signal init132_outs : std_logic_vector(31 downto 0);
  signal init132_outs_valid : std_logic;
  signal init132_outs_ready : std_logic;
  signal buffer9_outs_valid : std_logic;
  signal buffer9_outs_ready : std_logic;
  signal init133_outs_valid : std_logic;
  signal init133_outs_ready : std_logic;
  signal init134_outs_valid : std_logic;
  signal init134_outs_ready : std_logic;
  signal cond_br157_trueOut_valid : std_logic;
  signal cond_br157_trueOut_ready : std_logic;
  signal cond_br157_falseOut_valid : std_logic;
  signal cond_br157_falseOut_ready : std_logic;
  signal buffer226_outs : std_logic_vector(0 downto 0);
  signal buffer226_outs_valid : std_logic;
  signal buffer226_outs_ready : std_logic;
  signal cond_br158_trueOut_valid : std_logic;
  signal cond_br158_trueOut_ready : std_logic;
  signal cond_br158_falseOut_valid : std_logic;
  signal cond_br158_falseOut_ready : std_logic;
  signal buffer227_outs : std_logic_vector(0 downto 0);
  signal buffer227_outs_valid : std_logic;
  signal buffer227_outs_ready : std_logic;
  signal source15_outs_valid : std_logic;
  signal source15_outs_ready : std_logic;
  signal mux133_outs_valid : std_logic;
  signal mux133_outs_ready : std_logic;
  signal buffer228_outs : std_logic_vector(0 downto 0);
  signal buffer228_outs_valid : std_logic;
  signal buffer228_outs_ready : std_logic;
  signal source16_outs_valid : std_logic;
  signal source16_outs_ready : std_logic;
  signal mux134_outs_valid : std_logic;
  signal mux134_outs_ready : std_logic;
  signal buffer229_outs : std_logic_vector(0 downto 0);
  signal buffer229_outs_valid : std_logic;
  signal buffer229_outs_ready : std_logic;
  signal buffer103_outs_valid : std_logic;
  signal buffer103_outs_ready : std_logic;
  signal buffer104_outs_valid : std_logic;
  signal buffer104_outs_ready : std_logic;
  signal join4_outs_valid : std_logic;
  signal join4_outs_ready : std_logic;
  signal gate9_outs : std_logic_vector(31 downto 0);
  signal gate9_outs_valid : std_logic;
  signal gate9_outs_ready : std_logic;
  signal buffer230_outs : std_logic_vector(31 downto 0);
  signal buffer230_outs_valid : std_logic;
  signal buffer230_outs_ready : std_logic;
  signal trunci5_outs : std_logic_vector(6 downto 0);
  signal trunci5_outs_valid : std_logic;
  signal trunci5_outs_ready : std_logic;
  signal load3_addrOut : std_logic_vector(6 downto 0);
  signal load3_addrOut_valid : std_logic;
  signal load3_addrOut_ready : std_logic;
  signal load3_dataOut : std_logic_vector(31 downto 0);
  signal load3_dataOut_valid : std_logic;
  signal load3_dataOut_ready : std_logic;
  signal fork81_outs_0 : std_logic_vector(31 downto 0);
  signal fork81_outs_0_valid : std_logic;
  signal fork81_outs_0_ready : std_logic;
  signal fork81_outs_1 : std_logic_vector(31 downto 0);
  signal fork81_outs_1_valid : std_logic;
  signal fork81_outs_1_ready : std_logic;
  signal gate10_outs : std_logic_vector(31 downto 0);
  signal gate10_outs_valid : std_logic;
  signal gate10_outs_ready : std_logic;
  signal buffer231_outs : std_logic_vector(31 downto 0);
  signal buffer231_outs_valid : std_logic;
  signal buffer231_outs_ready : std_logic;
  signal fork82_outs_0 : std_logic_vector(31 downto 0);
  signal fork82_outs_0_valid : std_logic;
  signal fork82_outs_0_ready : std_logic;
  signal fork82_outs_1 : std_logic_vector(31 downto 0);
  signal fork82_outs_1_valid : std_logic;
  signal fork82_outs_1_ready : std_logic;
  signal cmpi13_result : std_logic_vector(0 downto 0);
  signal cmpi13_result_valid : std_logic;
  signal cmpi13_result_ready : std_logic;
  signal fork83_outs_0 : std_logic_vector(0 downto 0);
  signal fork83_outs_0_valid : std_logic;
  signal fork83_outs_0_ready : std_logic;
  signal fork83_outs_1 : std_logic_vector(0 downto 0);
  signal fork83_outs_1_valid : std_logic;
  signal fork83_outs_1_ready : std_logic;
  signal cmpi14_result : std_logic_vector(0 downto 0);
  signal cmpi14_result_valid : std_logic;
  signal cmpi14_result_ready : std_logic;
  signal buffer234_outs : std_logic_vector(31 downto 0);
  signal buffer234_outs_valid : std_logic;
  signal buffer234_outs_ready : std_logic;
  signal fork84_outs_0 : std_logic_vector(0 downto 0);
  signal fork84_outs_0_valid : std_logic;
  signal fork84_outs_0_ready : std_logic;
  signal fork84_outs_1 : std_logic_vector(0 downto 0);
  signal fork84_outs_1_valid : std_logic;
  signal fork84_outs_1_ready : std_logic;
  signal gate11_outs : std_logic_vector(31 downto 0);
  signal gate11_outs_valid : std_logic;
  signal gate11_outs_ready : std_logic;
  signal buffer235_outs : std_logic_vector(31 downto 0);
  signal buffer235_outs_valid : std_logic;
  signal buffer235_outs_ready : std_logic;
  signal fork85_outs_0 : std_logic_vector(31 downto 0);
  signal fork85_outs_0_valid : std_logic;
  signal fork85_outs_0_ready : std_logic;
  signal fork85_outs_1 : std_logic_vector(31 downto 0);
  signal fork85_outs_1_valid : std_logic;
  signal fork85_outs_1_ready : std_logic;
  signal cmpi15_result : std_logic_vector(0 downto 0);
  signal cmpi15_result_valid : std_logic;
  signal cmpi15_result_ready : std_logic;
  signal buffer236_outs : std_logic_vector(31 downto 0);
  signal buffer236_outs_valid : std_logic;
  signal buffer236_outs_ready : std_logic;
  signal fork86_outs_0 : std_logic_vector(0 downto 0);
  signal fork86_outs_0_valid : std_logic;
  signal fork86_outs_0_ready : std_logic;
  signal fork86_outs_1 : std_logic_vector(0 downto 0);
  signal fork86_outs_1_valid : std_logic;
  signal fork86_outs_1_ready : std_logic;
  signal cmpi16_result : std_logic_vector(0 downto 0);
  signal cmpi16_result_valid : std_logic;
  signal cmpi16_result_ready : std_logic;
  signal buffer238_outs : std_logic_vector(31 downto 0);
  signal buffer238_outs_valid : std_logic;
  signal buffer238_outs_ready : std_logic;
  signal fork87_outs_0 : std_logic_vector(0 downto 0);
  signal fork87_outs_0_valid : std_logic;
  signal fork87_outs_0_ready : std_logic;
  signal fork87_outs_1 : std_logic_vector(0 downto 0);
  signal fork87_outs_1_valid : std_logic;
  signal fork87_outs_1_ready : std_logic;
  signal gate12_outs : std_logic_vector(31 downto 0);
  signal gate12_outs_valid : std_logic;
  signal gate12_outs_ready : std_logic;
  signal buffer240_outs : std_logic_vector(31 downto 0);
  signal buffer240_outs_valid : std_logic;
  signal buffer240_outs_ready : std_logic;
  signal fork88_outs_0 : std_logic_vector(31 downto 0);
  signal fork88_outs_0_valid : std_logic;
  signal fork88_outs_0_ready : std_logic;
  signal fork88_outs_1 : std_logic_vector(31 downto 0);
  signal fork88_outs_1_valid : std_logic;
  signal fork88_outs_1_ready : std_logic;
  signal cmpi17_result : std_logic_vector(0 downto 0);
  signal cmpi17_result_valid : std_logic;
  signal cmpi17_result_ready : std_logic;
  signal fork89_outs_0 : std_logic_vector(0 downto 0);
  signal fork89_outs_0_valid : std_logic;
  signal fork89_outs_0_ready : std_logic;
  signal fork89_outs_1 : std_logic_vector(0 downto 0);
  signal fork89_outs_1_valid : std_logic;
  signal fork89_outs_1_ready : std_logic;
  signal cmpi18_result : std_logic_vector(0 downto 0);
  signal cmpi18_result_valid : std_logic;
  signal cmpi18_result_ready : std_logic;
  signal buffer243_outs : std_logic_vector(31 downto 0);
  signal buffer243_outs_valid : std_logic;
  signal buffer243_outs_ready : std_logic;
  signal fork90_outs_0 : std_logic_vector(0 downto 0);
  signal fork90_outs_0_valid : std_logic;
  signal fork90_outs_0_ready : std_logic;
  signal fork90_outs_1 : std_logic_vector(0 downto 0);
  signal fork90_outs_1_valid : std_logic;
  signal fork90_outs_1_ready : std_logic;
  signal buffer10_outs : std_logic_vector(7 downto 0);
  signal buffer10_outs_valid : std_logic;
  signal buffer10_outs_ready : std_logic;
  signal fork91_outs_0 : std_logic_vector(7 downto 0);
  signal fork91_outs_0_valid : std_logic;
  signal fork91_outs_0_ready : std_logic;
  signal fork91_outs_1 : std_logic_vector(7 downto 0);
  signal fork91_outs_1_valid : std_logic;
  signal fork91_outs_1_ready : std_logic;
  signal extsi44_outs : std_logic_vector(31 downto 0);
  signal extsi44_outs_valid : std_logic;
  signal extsi44_outs_ready : std_logic;
  signal buffer245_outs : std_logic_vector(7 downto 0);
  signal buffer245_outs_valid : std_logic;
  signal buffer245_outs_ready : std_logic;
  signal init135_outs : std_logic_vector(31 downto 0);
  signal init135_outs_valid : std_logic;
  signal init135_outs_ready : std_logic;
  signal buffer11_outs_valid : std_logic;
  signal buffer11_outs_ready : std_logic;
  signal init136_outs_valid : std_logic;
  signal init136_outs_ready : std_logic;
  signal fork92_outs_0_valid : std_logic;
  signal fork92_outs_0_ready : std_logic;
  signal fork92_outs_1_valid : std_logic;
  signal fork92_outs_1_ready : std_logic;
  signal init137_outs_valid : std_logic;
  signal init137_outs_ready : std_logic;
  signal cond_br159_trueOut_valid : std_logic;
  signal cond_br159_trueOut_ready : std_logic;
  signal cond_br159_falseOut_valid : std_logic;
  signal cond_br159_falseOut_ready : std_logic;
  signal cond_br160_trueOut_valid : std_logic;
  signal cond_br160_trueOut_ready : std_logic;
  signal cond_br160_falseOut_valid : std_logic;
  signal cond_br160_falseOut_ready : std_logic;
  signal buffer247_outs : std_logic_vector(0 downto 0);
  signal buffer247_outs_valid : std_logic;
  signal buffer247_outs_ready : std_logic;
  signal source17_outs_valid : std_logic;
  signal source17_outs_ready : std_logic;
  signal mux135_outs_valid : std_logic;
  signal mux135_outs_ready : std_logic;
  signal buffer248_outs : std_logic_vector(0 downto 0);
  signal buffer248_outs_valid : std_logic;
  signal buffer248_outs_ready : std_logic;
  signal source18_outs_valid : std_logic;
  signal source18_outs_ready : std_logic;
  signal mux136_outs_valid : std_logic;
  signal mux136_outs_ready : std_logic;
  signal buffer249_outs : std_logic_vector(0 downto 0);
  signal buffer249_outs_valid : std_logic;
  signal buffer249_outs_ready : std_logic;
  signal buffer105_outs_valid : std_logic;
  signal buffer105_outs_ready : std_logic;
  signal buffer106_outs_valid : std_logic;
  signal buffer106_outs_ready : std_logic;
  signal join5_outs_valid : std_logic;
  signal join5_outs_ready : std_logic;
  signal cond_br161_trueOut_valid : std_logic;
  signal cond_br161_trueOut_ready : std_logic;
  signal cond_br161_falseOut_valid : std_logic;
  signal cond_br161_falseOut_ready : std_logic;
  signal buffer250_outs : std_logic_vector(0 downto 0);
  signal buffer250_outs_valid : std_logic;
  signal buffer250_outs_ready : std_logic;
  signal cond_br162_trueOut_valid : std_logic;
  signal cond_br162_trueOut_ready : std_logic;
  signal cond_br162_falseOut_valid : std_logic;
  signal cond_br162_falseOut_ready : std_logic;
  signal buffer251_outs : std_logic_vector(0 downto 0);
  signal buffer251_outs_valid : std_logic;
  signal buffer251_outs_ready : std_logic;
  signal source19_outs_valid : std_logic;
  signal source19_outs_ready : std_logic;
  signal mux137_outs_valid : std_logic;
  signal mux137_outs_ready : std_logic;
  signal buffer252_outs : std_logic_vector(0 downto 0);
  signal buffer252_outs_valid : std_logic;
  signal buffer252_outs_ready : std_logic;
  signal source20_outs_valid : std_logic;
  signal source20_outs_ready : std_logic;
  signal mux138_outs_valid : std_logic;
  signal mux138_outs_ready : std_logic;
  signal buffer253_outs : std_logic_vector(0 downto 0);
  signal buffer253_outs_valid : std_logic;
  signal buffer253_outs_ready : std_logic;
  signal buffer107_outs_valid : std_logic;
  signal buffer107_outs_ready : std_logic;
  signal buffer108_outs_valid : std_logic;
  signal buffer108_outs_ready : std_logic;
  signal join6_outs_valid : std_logic;
  signal join6_outs_ready : std_logic;
  signal cond_br163_trueOut_valid : std_logic;
  signal cond_br163_trueOut_ready : std_logic;
  signal cond_br163_falseOut_valid : std_logic;
  signal cond_br163_falseOut_ready : std_logic;
  signal buffer254_outs : std_logic_vector(0 downto 0);
  signal buffer254_outs_valid : std_logic;
  signal buffer254_outs_ready : std_logic;
  signal cond_br164_trueOut_valid : std_logic;
  signal cond_br164_trueOut_ready : std_logic;
  signal cond_br164_falseOut_valid : std_logic;
  signal cond_br164_falseOut_ready : std_logic;
  signal buffer255_outs : std_logic_vector(0 downto 0);
  signal buffer255_outs_valid : std_logic;
  signal buffer255_outs_ready : std_logic;
  signal source21_outs_valid : std_logic;
  signal source21_outs_ready : std_logic;
  signal mux139_outs_valid : std_logic;
  signal mux139_outs_ready : std_logic;
  signal buffer256_outs : std_logic_vector(0 downto 0);
  signal buffer256_outs_valid : std_logic;
  signal buffer256_outs_ready : std_logic;
  signal source22_outs_valid : std_logic;
  signal source22_outs_ready : std_logic;
  signal mux140_outs_valid : std_logic;
  signal mux140_outs_ready : std_logic;
  signal buffer257_outs : std_logic_vector(0 downto 0);
  signal buffer257_outs_valid : std_logic;
  signal buffer257_outs_ready : std_logic;
  signal buffer109_outs_valid : std_logic;
  signal buffer109_outs_ready : std_logic;
  signal buffer110_outs_valid : std_logic;
  signal buffer110_outs_ready : std_logic;
  signal join7_outs_valid : std_logic;
  signal join7_outs_ready : std_logic;
  signal gate13_outs : std_logic_vector(31 downto 0);
  signal gate13_outs_valid : std_logic;
  signal gate13_outs_ready : std_logic;
  signal buffer258_outs : std_logic_vector(31 downto 0);
  signal buffer258_outs_valid : std_logic;
  signal buffer258_outs_ready : std_logic;
  signal buffer111_outs : std_logic_vector(31 downto 0);
  signal buffer111_outs_valid : std_logic;
  signal buffer111_outs_ready : std_logic;
  signal trunci6_outs : std_logic_vector(6 downto 0);
  signal trunci6_outs_valid : std_logic;
  signal trunci6_outs_ready : std_logic;
  signal store1_addrOut : std_logic_vector(6 downto 0);
  signal store1_addrOut_valid : std_logic;
  signal store1_addrOut_ready : std_logic;
  signal store1_dataToMem : std_logic_vector(31 downto 0);
  signal store1_dataToMem_valid : std_logic;
  signal store1_dataToMem_ready : std_logic;
  signal store1_doneOut_valid : std_logic;
  signal store1_doneOut_ready : std_logic;
  signal addi5_result : std_logic_vector(8 downto 0);
  signal addi5_result_valid : std_logic;
  signal addi5_result_ready : std_logic;
  signal buffer112_outs : std_logic_vector(8 downto 0);
  signal buffer112_outs_valid : std_logic;
  signal buffer112_outs_ready : std_logic;
  signal fork93_outs_0 : std_logic_vector(8 downto 0);
  signal fork93_outs_0_valid : std_logic;
  signal fork93_outs_0_ready : std_logic;
  signal fork93_outs_1 : std_logic_vector(8 downto 0);
  signal fork93_outs_1_valid : std_logic;
  signal fork93_outs_1_ready : std_logic;
  signal trunci7_outs : std_logic_vector(7 downto 0);
  signal trunci7_outs_valid : std_logic;
  signal trunci7_outs_ready : std_logic;
  signal buffer260_outs : std_logic_vector(8 downto 0);
  signal buffer260_outs_valid : std_logic;
  signal buffer260_outs_ready : std_logic;
  signal cmpi1_result : std_logic_vector(0 downto 0);
  signal cmpi1_result_valid : std_logic;
  signal cmpi1_result_ready : std_logic;
  signal buffer261_outs : std_logic_vector(8 downto 0);
  signal buffer261_outs_valid : std_logic;
  signal buffer261_outs_ready : std_logic;
  signal buffer113_outs : std_logic_vector(0 downto 0);
  signal buffer113_outs_valid : std_logic;
  signal buffer113_outs_ready : std_logic;
  signal fork94_outs_0 : std_logic_vector(0 downto 0);
  signal fork94_outs_0_valid : std_logic;
  signal fork94_outs_0_ready : std_logic;
  signal fork94_outs_1 : std_logic_vector(0 downto 0);
  signal fork94_outs_1_valid : std_logic;
  signal fork94_outs_1_ready : std_logic;
  signal fork94_outs_2 : std_logic_vector(0 downto 0);
  signal fork94_outs_2_valid : std_logic;
  signal fork94_outs_2_ready : std_logic;
  signal fork94_outs_3 : std_logic_vector(0 downto 0);
  signal fork94_outs_3_valid : std_logic;
  signal fork94_outs_3_ready : std_logic;
  signal fork94_outs_4 : std_logic_vector(0 downto 0);
  signal fork94_outs_4_valid : std_logic;
  signal fork94_outs_4_ready : std_logic;
  signal fork94_outs_5 : std_logic_vector(0 downto 0);
  signal fork94_outs_5_valid : std_logic;
  signal fork94_outs_5_ready : std_logic;
  signal fork94_outs_6 : std_logic_vector(0 downto 0);
  signal fork94_outs_6_valid : std_logic;
  signal fork94_outs_6_ready : std_logic;
  signal fork94_outs_7 : std_logic_vector(0 downto 0);
  signal fork94_outs_7_valid : std_logic;
  signal fork94_outs_7_ready : std_logic;
  signal fork94_outs_8 : std_logic_vector(0 downto 0);
  signal fork94_outs_8_valid : std_logic;
  signal fork94_outs_8_ready : std_logic;
  signal fork94_outs_9 : std_logic_vector(0 downto 0);
  signal fork94_outs_9_valid : std_logic;
  signal fork94_outs_9_ready : std_logic;
  signal fork94_outs_10 : std_logic_vector(0 downto 0);
  signal fork94_outs_10_valid : std_logic;
  signal fork94_outs_10_ready : std_logic;
  signal fork94_outs_11 : std_logic_vector(0 downto 0);
  signal fork94_outs_11_valid : std_logic;
  signal fork94_outs_11_ready : std_logic;
  signal fork94_outs_12 : std_logic_vector(0 downto 0);
  signal fork94_outs_12_valid : std_logic;
  signal fork94_outs_12_ready : std_logic;
  signal fork94_outs_13 : std_logic_vector(0 downto 0);
  signal fork94_outs_13_valid : std_logic;
  signal fork94_outs_13_ready : std_logic;
  signal fork94_outs_14 : std_logic_vector(0 downto 0);
  signal fork94_outs_14_valid : std_logic;
  signal fork94_outs_14_ready : std_logic;
  signal fork94_outs_15 : std_logic_vector(0 downto 0);
  signal fork94_outs_15_valid : std_logic;
  signal fork94_outs_15_ready : std_logic;
  signal fork94_outs_16 : std_logic_vector(0 downto 0);
  signal fork94_outs_16_valid : std_logic;
  signal fork94_outs_16_ready : std_logic;
  signal fork94_outs_17 : std_logic_vector(0 downto 0);
  signal fork94_outs_17_valid : std_logic;
  signal fork94_outs_17_ready : std_logic;
  signal fork94_outs_18 : std_logic_vector(0 downto 0);
  signal fork94_outs_18_valid : std_logic;
  signal fork94_outs_18_ready : std_logic;
  signal fork94_outs_19 : std_logic_vector(0 downto 0);
  signal fork94_outs_19_valid : std_logic;
  signal fork94_outs_19_ready : std_logic;
  signal fork94_outs_20 : std_logic_vector(0 downto 0);
  signal fork94_outs_20_valid : std_logic;
  signal fork94_outs_20_ready : std_logic;
  signal fork94_outs_21 : std_logic_vector(0 downto 0);
  signal fork94_outs_21_valid : std_logic;
  signal fork94_outs_21_ready : std_logic;
  signal fork94_outs_22 : std_logic_vector(0 downto 0);
  signal fork94_outs_22_valid : std_logic;
  signal fork94_outs_22_ready : std_logic;
  signal fork94_outs_23 : std_logic_vector(0 downto 0);
  signal fork94_outs_23_valid : std_logic;
  signal fork94_outs_23_ready : std_logic;
  signal fork94_outs_24 : std_logic_vector(0 downto 0);
  signal fork94_outs_24_valid : std_logic;
  signal fork94_outs_24_ready : std_logic;
  signal fork94_outs_25 : std_logic_vector(0 downto 0);
  signal fork94_outs_25_valid : std_logic;
  signal fork94_outs_25_ready : std_logic;
  signal fork94_outs_26 : std_logic_vector(0 downto 0);
  signal fork94_outs_26_valid : std_logic;
  signal fork94_outs_26_ready : std_logic;
  signal fork94_outs_27 : std_logic_vector(0 downto 0);
  signal fork94_outs_27_valid : std_logic;
  signal fork94_outs_27_ready : std_logic;
  signal fork94_outs_28 : std_logic_vector(0 downto 0);
  signal fork94_outs_28_valid : std_logic;
  signal fork94_outs_28_ready : std_logic;
  signal cond_br7_trueOut : std_logic_vector(7 downto 0);
  signal cond_br7_trueOut_valid : std_logic;
  signal cond_br7_trueOut_ready : std_logic;
  signal cond_br7_falseOut : std_logic_vector(7 downto 0);
  signal cond_br7_falseOut_valid : std_logic;
  signal cond_br7_falseOut_ready : std_logic;
  signal buffer100_outs : std_logic_vector(2 downto 0);
  signal buffer100_outs_valid : std_logic;
  signal buffer100_outs_ready : std_logic;
  signal buffer101_outs : std_logic_vector(2 downto 0);
  signal buffer101_outs_valid : std_logic;
  signal buffer101_outs_ready : std_logic;
  signal cond_br8_trueOut : std_logic_vector(2 downto 0);
  signal cond_br8_trueOut_valid : std_logic;
  signal cond_br8_trueOut_ready : std_logic;
  signal cond_br8_falseOut : std_logic_vector(2 downto 0);
  signal cond_br8_falseOut_valid : std_logic;
  signal cond_br8_falseOut_ready : std_logic;
  signal buffer102_outs_valid : std_logic;
  signal buffer102_outs_ready : std_logic;
  signal cond_br9_trueOut_valid : std_logic;
  signal cond_br9_trueOut_ready : std_logic;
  signal cond_br9_falseOut_valid : std_logic;
  signal cond_br9_falseOut_ready : std_logic;
  signal buffer264_outs : std_logic_vector(0 downto 0);
  signal buffer264_outs_valid : std_logic;
  signal buffer264_outs_ready : std_logic;
  signal cond_br259_trueOut : std_logic_vector(31 downto 0);
  signal cond_br259_trueOut_valid : std_logic;
  signal cond_br259_trueOut_ready : std_logic;
  signal cond_br259_falseOut : std_logic_vector(31 downto 0);
  signal cond_br259_falseOut_valid : std_logic;
  signal cond_br259_falseOut_ready : std_logic;
  signal fork95_outs_0 : std_logic_vector(31 downto 0);
  signal fork95_outs_0_valid : std_logic;
  signal fork95_outs_0_ready : std_logic;
  signal fork95_outs_1 : std_logic_vector(31 downto 0);
  signal fork95_outs_1_valid : std_logic;
  signal fork95_outs_1_ready : std_logic;
  signal fork95_outs_2 : std_logic_vector(31 downto 0);
  signal fork95_outs_2_valid : std_logic;
  signal fork95_outs_2_ready : std_logic;
  signal cond_br260_trueOut : std_logic_vector(7 downto 0);
  signal cond_br260_trueOut_valid : std_logic;
  signal cond_br260_trueOut_ready : std_logic;
  signal cond_br260_falseOut : std_logic_vector(7 downto 0);
  signal cond_br260_falseOut_valid : std_logic;
  signal cond_br260_falseOut_ready : std_logic;
  signal fork96_outs_0 : std_logic_vector(7 downto 0);
  signal fork96_outs_0_valid : std_logic;
  signal fork96_outs_0_ready : std_logic;
  signal fork96_outs_1 : std_logic_vector(7 downto 0);
  signal fork96_outs_1_valid : std_logic;
  signal fork96_outs_1_ready : std_logic;
  signal fork96_outs_2 : std_logic_vector(7 downto 0);
  signal fork96_outs_2_valid : std_logic;
  signal fork96_outs_2_ready : std_logic;
  signal extsi45_outs : std_logic_vector(10 downto 0);
  signal extsi45_outs_valid : std_logic;
  signal extsi45_outs_ready : std_logic;
  signal extsi46_outs : std_logic_vector(10 downto 0);
  signal extsi46_outs_valid : std_logic;
  signal extsi46_outs_ready : std_logic;
  signal extsi47_outs : std_logic_vector(10 downto 0);
  signal extsi47_outs_valid : std_logic;
  signal extsi47_outs_ready : std_logic;
  signal cond_br261_trueOut : std_logic_vector(7 downto 0);
  signal cond_br261_trueOut_valid : std_logic;
  signal cond_br261_trueOut_ready : std_logic;
  signal cond_br261_falseOut : std_logic_vector(7 downto 0);
  signal cond_br261_falseOut_valid : std_logic;
  signal cond_br261_falseOut_ready : std_logic;
  signal extsi48_outs : std_logic_vector(10 downto 0);
  signal extsi48_outs_valid : std_logic;
  signal extsi48_outs_ready : std_logic;
  signal cond_br262_trueOut : std_logic_vector(31 downto 0);
  signal cond_br262_trueOut_valid : std_logic;
  signal cond_br262_trueOut_ready : std_logic;
  signal cond_br262_falseOut : std_logic_vector(31 downto 0);
  signal cond_br262_falseOut_valid : std_logic;
  signal cond_br262_falseOut_ready : std_logic;
  signal cond_br263_trueOut_valid : std_logic;
  signal cond_br263_trueOut_ready : std_logic;
  signal cond_br263_falseOut_valid : std_logic;
  signal cond_br263_falseOut_ready : std_logic;
  signal buffer272_outs : std_logic_vector(0 downto 0);
  signal buffer272_outs_valid : std_logic;
  signal buffer272_outs_ready : std_logic;
  signal extsi49_outs : std_logic_vector(3 downto 0);
  signal extsi49_outs_valid : std_logic;
  signal extsi49_outs_ready : std_logic;
  signal source5_outs_valid : std_logic;
  signal source5_outs_ready : std_logic;
  signal constant29_outs : std_logic_vector(2 downto 0);
  signal constant29_outs_valid : std_logic;
  signal constant29_outs_ready : std_logic;
  signal extsi50_outs : std_logic_vector(3 downto 0);
  signal extsi50_outs_valid : std_logic;
  signal extsi50_outs_ready : std_logic;
  signal source6_outs_valid : std_logic;
  signal source6_outs_ready : std_logic;
  signal constant30_outs : std_logic_vector(1 downto 0);
  signal constant30_outs_valid : std_logic;
  signal constant30_outs_ready : std_logic;
  signal extsi51_outs : std_logic_vector(3 downto 0);
  signal extsi51_outs_valid : std_logic;
  signal extsi51_outs_ready : std_logic;
  signal addi6_result : std_logic_vector(3 downto 0);
  signal addi6_result_valid : std_logic;
  signal addi6_result_ready : std_logic;
  signal buffer114_outs : std_logic_vector(3 downto 0);
  signal buffer114_outs_valid : std_logic;
  signal buffer114_outs_ready : std_logic;
  signal fork97_outs_0 : std_logic_vector(3 downto 0);
  signal fork97_outs_0_valid : std_logic;
  signal fork97_outs_0_ready : std_logic;
  signal fork97_outs_1 : std_logic_vector(3 downto 0);
  signal fork97_outs_1_valid : std_logic;
  signal fork97_outs_1_ready : std_logic;
  signal trunci8_outs : std_logic_vector(2 downto 0);
  signal trunci8_outs_valid : std_logic;
  signal trunci8_outs_ready : std_logic;
  signal cmpi2_result : std_logic_vector(0 downto 0);
  signal cmpi2_result_valid : std_logic;
  signal cmpi2_result_ready : std_logic;
  signal buffer115_outs : std_logic_vector(0 downto 0);
  signal buffer115_outs_valid : std_logic;
  signal buffer115_outs_ready : std_logic;
  signal fork98_outs_0 : std_logic_vector(0 downto 0);
  signal fork98_outs_0_valid : std_logic;
  signal fork98_outs_0_ready : std_logic;
  signal fork98_outs_1 : std_logic_vector(0 downto 0);
  signal fork98_outs_1_valid : std_logic;
  signal fork98_outs_1_ready : std_logic;
  signal fork98_outs_2 : std_logic_vector(0 downto 0);
  signal fork98_outs_2_valid : std_logic;
  signal fork98_outs_2_ready : std_logic;
  signal fork98_outs_3 : std_logic_vector(0 downto 0);
  signal fork98_outs_3_valid : std_logic;
  signal fork98_outs_3_ready : std_logic;
  signal fork98_outs_4 : std_logic_vector(0 downto 0);
  signal fork98_outs_4_valid : std_logic;
  signal fork98_outs_4_ready : std_logic;
  signal fork98_outs_5 : std_logic_vector(0 downto 0);
  signal fork98_outs_5_valid : std_logic;
  signal fork98_outs_5_ready : std_logic;
  signal fork98_outs_6 : std_logic_vector(0 downto 0);
  signal fork98_outs_6_valid : std_logic;
  signal fork98_outs_6_ready : std_logic;
  signal fork98_outs_7 : std_logic_vector(0 downto 0);
  signal fork98_outs_7_valid : std_logic;
  signal fork98_outs_7_ready : std_logic;
  signal cond_br10_trueOut : std_logic_vector(2 downto 0);
  signal cond_br10_trueOut_valid : std_logic;
  signal cond_br10_trueOut_ready : std_logic;
  signal cond_br10_falseOut : std_logic_vector(2 downto 0);
  signal cond_br10_falseOut_valid : std_logic;
  signal cond_br10_falseOut_ready : std_logic;
  signal cond_br11_trueOut_valid : std_logic;
  signal cond_br11_trueOut_ready : std_logic;
  signal cond_br11_falseOut_valid : std_logic;
  signal cond_br11_falseOut_ready : std_logic;
  signal buffer276_outs : std_logic_vector(0 downto 0);
  signal buffer276_outs_valid : std_logic;
  signal buffer276_outs_ready : std_logic;
  signal fork99_outs_0_valid : std_logic;
  signal fork99_outs_0_ready : std_logic;
  signal fork99_outs_1_valid : std_logic;
  signal fork99_outs_1_ready : std_logic;

begin

  A_end_valid <= mem_controller1_memEnd_valid;
  mem_controller1_memEnd_ready <= A_end_ready;
  B_end_valid <= mem_controller0_memEnd_valid;
  mem_controller0_memEnd_ready <= B_end_ready;
  end_valid <= fork0_outs_2_valid;
  fork0_outs_2_ready <= end_ready;
  A_loadEn <= mem_controller1_loadEn;
  A_loadAddr <= mem_controller1_loadAddr;
  A_storeEn <= mem_controller1_storeEn;
  A_storeAddr <= mem_controller1_storeAddr;
  A_storeData <= mem_controller1_storeData;
  B_loadEn <= mem_controller0_loadEn;
  B_loadAddr <= mem_controller0_loadAddr;
  B_storeEn <= mem_controller0_storeEn;
  B_storeAddr <= mem_controller0_storeAddr;
  B_storeData <= mem_controller0_storeData;

  fork0 : entity work.fork_dataless(arch) generic map(5)
    port map(
      ins_valid => start_valid,
      ins_ready => start_ready,
      clk => clk,
      rst => rst,
      outs_valid(0) => fork0_outs_0_valid,
      outs_valid(1) => fork0_outs_1_valid,
      outs_valid(2) => fork0_outs_2_valid,
      outs_valid(3) => fork0_outs_3_valid,
      outs_valid(4) => fork0_outs_4_valid,
      outs_ready(0) => fork0_outs_0_ready,
      outs_ready(1) => fork0_outs_1_ready,
      outs_ready(2) => fork0_outs_2_ready,
      outs_ready(3) => fork0_outs_3_ready,
      outs_ready(4) => fork0_outs_4_ready
    );

  mem_controller0 : entity work.mem_controller(arch) generic map(1, 1, 1, 32, 7)
    port map(
      loadData => B_loadData,
      memStart_valid => B_start_valid,
      memStart_ready => B_start_ready,
      ctrl(0) => extsi11_outs,
      ctrl_valid(0) => extsi11_outs_valid,
      ctrl_ready(0) => extsi11_outs_ready,
      stAddr(0) => store0_addrOut,
      stAddr_valid(0) => store0_addrOut_valid,
      stAddr_ready(0) => store0_addrOut_ready,
      stData(0) => store0_dataToMem,
      stData_valid(0) => store0_dataToMem_valid,
      stData_ready(0) => store0_dataToMem_ready,
      ldAddr(0) => load3_addrOut,
      ldAddr_valid(0) => load3_addrOut_valid,
      ldAddr_ready(0) => load3_addrOut_ready,
      ctrlEnd_valid => fork99_outs_1_valid,
      ctrlEnd_ready => fork99_outs_1_ready,
      clk => clk,
      rst => rst,
      stDone_valid(0) => mem_controller0_stDone_0_valid,
      stDone_ready(0) => mem_controller0_stDone_0_ready,
      ldData(0) => mem_controller0_ldData_0,
      ldData_valid(0) => mem_controller0_ldData_0_valid,
      ldData_ready(0) => mem_controller0_ldData_0_ready,
      memEnd_valid => mem_controller0_memEnd_valid,
      memEnd_ready => mem_controller0_memEnd_ready,
      loadEn => mem_controller0_loadEn,
      loadAddr => mem_controller0_loadAddr,
      storeEn => mem_controller0_storeEn,
      storeAddr => mem_controller0_storeAddr,
      storeData => mem_controller0_storeData
    );

  mem_controller1 : entity work.mem_controller(arch) generic map(1, 3, 1, 32, 7)
    port map(
      loadData => A_loadData,
      memStart_valid => A_start_valid,
      memStart_ready => A_start_ready,
      ldAddr(0) => load0_addrOut,
      ldAddr(1) => load1_addrOut,
      ldAddr(2) => load2_addrOut,
      ldAddr_valid(0) => load0_addrOut_valid,
      ldAddr_valid(1) => load1_addrOut_valid,
      ldAddr_valid(2) => load2_addrOut_valid,
      ldAddr_ready(0) => load0_addrOut_ready,
      ldAddr_ready(1) => load1_addrOut_ready,
      ldAddr_ready(2) => load2_addrOut_ready,
      ctrl(0) => extsi14_outs,
      ctrl_valid(0) => extsi14_outs_valid,
      ctrl_ready(0) => extsi14_outs_ready,
      stAddr(0) => store1_addrOut,
      stAddr_valid(0) => store1_addrOut_valid,
      stAddr_ready(0) => store1_addrOut_ready,
      stData(0) => store1_dataToMem,
      stData_valid(0) => store1_dataToMem_valid,
      stData_ready(0) => store1_dataToMem_ready,
      ctrlEnd_valid => fork99_outs_0_valid,
      ctrlEnd_ready => fork99_outs_0_ready,
      clk => clk,
      rst => rst,
      ldData(0) => mem_controller1_ldData_0,
      ldData(1) => mem_controller1_ldData_1,
      ldData(2) => mem_controller1_ldData_2,
      ldData_valid(0) => mem_controller1_ldData_0_valid,
      ldData_valid(1) => mem_controller1_ldData_1_valid,
      ldData_valid(2) => mem_controller1_ldData_2_valid,
      ldData_ready(0) => mem_controller1_ldData_0_ready,
      ldData_ready(1) => mem_controller1_ldData_1_ready,
      ldData_ready(2) => mem_controller1_ldData_2_ready,
      stDone_valid(0) => mem_controller1_stDone_0_valid,
      stDone_ready(0) => mem_controller1_stDone_0_ready,
      memEnd_valid => mem_controller1_memEnd_valid,
      memEnd_ready => mem_controller1_memEnd_ready,
      loadEn => mem_controller1_loadEn,
      loadAddr => mem_controller1_loadAddr,
      storeEn => mem_controller1_storeEn,
      storeAddr => mem_controller1_storeAddr,
      storeData => mem_controller1_storeData
    );

  constant1 : entity work.handshake_constant_0(arch) generic map(11)
    port map(
      ctrl_valid => fork0_outs_1_valid,
      ctrl_ready => fork0_outs_1_ready,
      clk => clk,
      rst => rst,
      outs => constant1_outs,
      outs_valid => constant1_outs_valid,
      outs_ready => constant1_outs_ready
    );

  fork1 : entity work.handshake_fork(arch) generic map(8, 11)
    port map(
      ins => constant1_outs,
      ins_valid => constant1_outs_valid,
      ins_ready => constant1_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork1_outs_0,
      outs(1) => fork1_outs_1,
      outs(2) => fork1_outs_2,
      outs(3) => fork1_outs_3,
      outs(4) => fork1_outs_4,
      outs(5) => fork1_outs_5,
      outs(6) => fork1_outs_6,
      outs(7) => fork1_outs_7,
      outs_valid(0) => fork1_outs_0_valid,
      outs_valid(1) => fork1_outs_1_valid,
      outs_valid(2) => fork1_outs_2_valid,
      outs_valid(3) => fork1_outs_3_valid,
      outs_valid(4) => fork1_outs_4_valid,
      outs_valid(5) => fork1_outs_5_valid,
      outs_valid(6) => fork1_outs_6_valid,
      outs_valid(7) => fork1_outs_7_valid,
      outs_ready(0) => fork1_outs_0_ready,
      outs_ready(1) => fork1_outs_1_ready,
      outs_ready(2) => fork1_outs_2_ready,
      outs_ready(3) => fork1_outs_3_ready,
      outs_ready(4) => fork1_outs_4_ready,
      outs_ready(5) => fork1_outs_5_ready,
      outs_ready(6) => fork1_outs_6_ready,
      outs_ready(7) => fork1_outs_7_ready
    );

  extsi0 : entity work.extsi(arch) generic map(11, 32)
    port map(
      ins => fork1_outs_4,
      ins_valid => fork1_outs_4_valid,
      ins_ready => fork1_outs_4_ready,
      clk => clk,
      rst => rst,
      outs => extsi0_outs,
      outs_valid => extsi0_outs_valid,
      outs_ready => extsi0_outs_ready
    );

  extsi1 : entity work.extsi(arch) generic map(11, 32)
    port map(
      ins => fork1_outs_5,
      ins_valid => fork1_outs_5_valid,
      ins_ready => fork1_outs_5_ready,
      clk => clk,
      rst => rst,
      outs => extsi1_outs,
      outs_valid => extsi1_outs_valid,
      outs_ready => extsi1_outs_ready
    );

  extsi5 : entity work.extsi(arch) generic map(11, 32)
    port map(
      ins => fork1_outs_6,
      ins_valid => fork1_outs_6_valid,
      ins_ready => fork1_outs_6_ready,
      clk => clk,
      rst => rst,
      outs => extsi5_outs,
      outs_valid => extsi5_outs_valid,
      outs_ready => extsi5_outs_ready
    );

  extsi6 : entity work.extsi(arch) generic map(11, 32)
    port map(
      ins => fork1_outs_7,
      ins_valid => fork1_outs_7_valid,
      ins_ready => fork1_outs_7_ready,
      clk => clk,
      rst => rst,
      outs => extsi6_outs,
      outs_valid => extsi6_outs_valid,
      outs_ready => extsi6_outs_ready
    );

  constant2 : entity work.handshake_constant_1(arch) generic map(1)
    port map(
      ctrl_valid => fork0_outs_0_valid,
      ctrl_ready => fork0_outs_0_ready,
      clk => clk,
      rst => rst,
      outs => constant2_outs,
      outs_valid => constant2_outs_valid,
      outs_ready => constant2_outs_ready
    );

  extsi21 : entity work.extsi(arch) generic map(1, 3)
    port map(
      ins => constant2_outs,
      ins_valid => constant2_outs_valid,
      ins_ready => constant2_outs_ready,
      clk => clk,
      rst => rst,
      outs => extsi21_outs,
      outs_valid => extsi21_outs_valid,
      outs_ready => extsi21_outs_ready
    );

  mux6 : entity work.mux(arch) generic map(2, 32, 1)
    port map(
      index => fork2_outs_4,
      index_valid => fork2_outs_4_valid,
      index_ready => fork2_outs_4_ready,
      ins(0) => extsi0_outs,
      ins(1) => fork95_outs_0,
      ins_valid(0) => extsi0_outs_valid,
      ins_valid(1) => fork95_outs_0_valid,
      ins_ready(0) => extsi0_outs_ready,
      ins_ready(1) => fork95_outs_0_ready,
      clk => clk,
      rst => rst,
      outs => mux6_outs,
      outs_valid => mux6_outs_valid,
      outs_ready => mux6_outs_ready
    );

  mux7 : entity work.mux(arch) generic map(2, 32, 1)
    port map(
      index => fork2_outs_5,
      index_valid => fork2_outs_5_valid,
      index_ready => fork2_outs_5_ready,
      ins(0) => extsi1_outs,
      ins(1) => fork95_outs_1,
      ins_valid(0) => extsi1_outs_valid,
      ins_valid(1) => fork95_outs_1_valid,
      ins_ready(0) => extsi1_outs_ready,
      ins_ready(1) => fork95_outs_1_ready,
      clk => clk,
      rst => rst,
      outs => mux7_outs,
      outs_valid => mux7_outs_valid,
      outs_ready => mux7_outs_ready
    );

  mux9 : entity work.mux(arch) generic map(2, 11, 1)
    port map(
      index => fork2_outs_0,
      index_valid => fork2_outs_0_valid,
      index_ready => fork2_outs_0_ready,
      ins(0) => fork1_outs_0,
      ins(1) => extsi45_outs,
      ins_valid(0) => fork1_outs_0_valid,
      ins_valid(1) => extsi45_outs_valid,
      ins_ready(0) => fork1_outs_0_ready,
      ins_ready(1) => extsi45_outs_ready,
      clk => clk,
      rst => rst,
      outs => mux9_outs,
      outs_valid => mux9_outs_valid,
      outs_ready => mux9_outs_ready
    );

  mux10 : entity work.mux(arch) generic map(2, 11, 1)
    port map(
      index => fork2_outs_1,
      index_valid => fork2_outs_1_valid,
      index_ready => fork2_outs_1_ready,
      ins(0) => fork1_outs_1,
      ins(1) => extsi46_outs,
      ins_valid(0) => fork1_outs_1_valid,
      ins_valid(1) => extsi46_outs_valid,
      ins_ready(0) => fork1_outs_1_ready,
      ins_ready(1) => extsi46_outs_ready,
      clk => clk,
      rst => rst,
      outs => mux10_outs,
      outs_valid => mux10_outs_valid,
      outs_ready => mux10_outs_ready
    );

  mux19 : entity work.mux(arch) generic map(2, 11, 1)
    port map(
      index => fork2_outs_2,
      index_valid => fork2_outs_2_valid,
      index_ready => fork2_outs_2_ready,
      ins(0) => fork1_outs_2,
      ins(1) => extsi48_outs,
      ins_valid(0) => fork1_outs_2_valid,
      ins_valid(1) => extsi48_outs_valid,
      ins_ready(0) => fork1_outs_2_ready,
      ins_ready(1) => extsi48_outs_ready,
      clk => clk,
      rst => rst,
      outs => mux19_outs,
      outs_valid => mux19_outs_valid,
      outs_ready => mux19_outs_ready
    );

  mux21 : entity work.mux(arch) generic map(2, 32, 1)
    port map(
      index => fork2_outs_6,
      index_valid => fork2_outs_6_valid,
      index_ready => fork2_outs_6_ready,
      ins(0) => extsi5_outs,
      ins(1) => fork95_outs_2,
      ins_valid(0) => extsi5_outs_valid,
      ins_valid(1) => fork95_outs_2_valid,
      ins_ready(0) => extsi5_outs_ready,
      ins_ready(1) => fork95_outs_2_ready,
      clk => clk,
      rst => rst,
      outs => mux21_outs,
      outs_valid => mux21_outs_valid,
      outs_ready => mux21_outs_ready
    );

  mux23 : entity work.mux(arch) generic map(2, 32, 1)
    port map(
      index => fork2_outs_7,
      index_valid => fork2_outs_7_valid,
      index_ready => fork2_outs_7_ready,
      ins(0) => extsi6_outs,
      ins(1) => cond_br262_trueOut,
      ins_valid(0) => extsi6_outs_valid,
      ins_valid(1) => cond_br262_trueOut_valid,
      ins_ready(0) => extsi6_outs_ready,
      ins_ready(1) => cond_br262_trueOut_ready,
      clk => clk,
      rst => rst,
      outs => mux23_outs,
      outs_valid => mux23_outs_valid,
      outs_ready => mux23_outs_ready
    );

  mux28 : entity work.mux(arch) generic map(2, 11, 1)
    port map(
      index => fork2_outs_3,
      index_valid => fork2_outs_3_valid,
      index_ready => fork2_outs_3_ready,
      ins(0) => fork1_outs_3,
      ins(1) => extsi47_outs,
      ins_valid(0) => fork1_outs_3_valid,
      ins_valid(1) => extsi47_outs_valid,
      ins_ready(0) => fork1_outs_3_ready,
      ins_ready(1) => extsi47_outs_ready,
      clk => clk,
      rst => rst,
      outs => mux28_outs,
      outs_valid => mux28_outs_valid,
      outs_ready => mux28_outs_ready
    );

  mux37 : entity work.mux_dataless(arch) generic map(2, 1)
    port map(
      index => fork2_outs_8,
      index_valid => fork2_outs_8_valid,
      index_ready => fork2_outs_8_ready,
      ins_valid(0) => fork0_outs_3_valid,
      ins_valid(1) => cond_br263_trueOut_valid,
      ins_ready(0) => fork0_outs_3_ready,
      ins_ready(1) => cond_br263_trueOut_ready,
      clk => clk,
      rst => rst,
      outs_valid => mux37_outs_valid,
      outs_ready => mux37_outs_ready
    );

  init0 : entity work.tehb_init(arch) generic map(1, 0)
    port map(
      ins => fork98_outs_4,
      ins_valid => fork98_outs_4_valid,
      ins_ready => fork98_outs_4_ready,
      clk => clk,
      rst => rst,
      outs => init0_outs,
      outs_valid => init0_outs_valid,
      outs_ready => init0_outs_ready
    );

  fork2 : entity work.handshake_fork(arch) generic map(9, 1)
    port map(
      ins => init0_outs,
      ins_valid => init0_outs_valid,
      ins_ready => init0_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork2_outs_0,
      outs(1) => fork2_outs_1,
      outs(2) => fork2_outs_2,
      outs(3) => fork2_outs_3,
      outs(4) => fork2_outs_4,
      outs(5) => fork2_outs_5,
      outs(6) => fork2_outs_6,
      outs(7) => fork2_outs_7,
      outs(8) => fork2_outs_8,
      outs_valid(0) => fork2_outs_0_valid,
      outs_valid(1) => fork2_outs_1_valid,
      outs_valid(2) => fork2_outs_2_valid,
      outs_valid(3) => fork2_outs_3_valid,
      outs_valid(4) => fork2_outs_4_valid,
      outs_valid(5) => fork2_outs_5_valid,
      outs_valid(6) => fork2_outs_6_valid,
      outs_valid(7) => fork2_outs_7_valid,
      outs_valid(8) => fork2_outs_8_valid,
      outs_ready(0) => fork2_outs_0_ready,
      outs_ready(1) => fork2_outs_1_ready,
      outs_ready(2) => fork2_outs_2_ready,
      outs_ready(3) => fork2_outs_3_ready,
      outs_ready(4) => fork2_outs_4_ready,
      outs_ready(5) => fork2_outs_5_ready,
      outs_ready(6) => fork2_outs_6_ready,
      outs_ready(7) => fork2_outs_7_ready,
      outs_ready(8) => fork2_outs_8_ready
    );

  mux0 : entity work.mux(arch) generic map(2, 3, 1)
    port map(
      index => control_merge0_index,
      index_valid => control_merge0_index_valid,
      index_ready => control_merge0_index_ready,
      ins(0) => extsi21_outs,
      ins(1) => cond_br10_trueOut,
      ins_valid(0) => extsi21_outs_valid,
      ins_valid(1) => cond_br10_trueOut_valid,
      ins_ready(0) => extsi21_outs_ready,
      ins_ready(1) => cond_br10_trueOut_ready,
      clk => clk,
      rst => rst,
      outs => mux0_outs,
      outs_valid => mux0_outs_valid,
      outs_ready => mux0_outs_ready
    );

  control_merge0 : entity work.control_merge_dataless(arch) generic map(2, 1)
    port map(
      ins_valid(0) => fork0_outs_4_valid,
      ins_valid(1) => cond_br11_trueOut_valid,
      ins_ready(0) => fork0_outs_4_ready,
      ins_ready(1) => cond_br11_trueOut_ready,
      clk => clk,
      rst => rst,
      outs_valid => control_merge0_outs_valid,
      outs_ready => control_merge0_outs_ready,
      index => control_merge0_index,
      index_valid => control_merge0_index_valid,
      index_ready => control_merge0_index_ready
    );

  fork3 : entity work.fork_dataless(arch) generic map(2)
    port map(
      ins_valid => control_merge0_outs_valid,
      ins_ready => control_merge0_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid(0) => fork3_outs_0_valid,
      outs_valid(1) => fork3_outs_1_valid,
      outs_ready(0) => fork3_outs_0_ready,
      outs_ready(1) => fork3_outs_1_ready
    );

  constant5 : entity work.handshake_constant_2(arch) generic map(2)
    port map(
      ctrl_valid => fork3_outs_0_valid,
      ctrl_ready => fork3_outs_0_ready,
      clk => clk,
      rst => rst,
      outs => constant5_outs,
      outs_valid => constant5_outs_valid,
      outs_ready => constant5_outs_ready
    );

  extsi20 : entity work.extsi(arch) generic map(2, 8)
    port map(
      ins => constant5_outs,
      ins_valid => constant5_outs_valid,
      ins_ready => constant5_outs_ready,
      clk => clk,
      rst => rst,
      outs => extsi20_outs,
      outs_valid => extsi20_outs_valid,
      outs_ready => extsi20_outs_ready
    );

  buffer13 : entity work.tehb(arch) generic map(3)
    port map(
      ins => mux0_outs,
      ins_valid => mux0_outs_valid,
      ins_ready => mux0_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer13_outs,
      outs_valid => buffer13_outs_valid,
      outs_ready => buffer13_outs_ready
    );

  cond_br205 : entity work.cond_br(arch) generic map(32)
    port map(
      condition => fork51_outs_31,
      condition_valid => fork51_outs_31_valid,
      condition_ready => fork51_outs_31_ready,
      data => fork11_outs_1,
      data_valid => fork11_outs_1_valid,
      data_ready => fork11_outs_1_ready,
      clk => clk,
      rst => rst,
      trueOut => cond_br205_trueOut,
      trueOut_valid => cond_br205_trueOut_valid,
      trueOut_ready => cond_br205_trueOut_ready,
      falseOut => cond_br205_falseOut,
      falseOut_valid => cond_br205_falseOut_valid,
      falseOut_ready => cond_br205_falseOut_ready
    );

  sink0 : entity work.sink(arch) generic map(32)
    port map(
      ins => cond_br205_falseOut,
      ins_valid => cond_br205_falseOut_valid,
      ins_ready => cond_br205_falseOut_ready,
      clk => clk,
      rst => rst
    );

  cond_br206 : entity work.cond_br_dataless(arch)
    port map(
      condition => fork51_outs_30,
      condition_valid => fork51_outs_30_valid,
      condition_ready => fork51_outs_30_ready,
      data_valid => fork29_outs_1_valid,
      data_ready => fork29_outs_1_ready,
      clk => clk,
      rst => rst,
      trueOut_valid => cond_br206_trueOut_valid,
      trueOut_ready => cond_br206_trueOut_ready,
      falseOut_valid => cond_br206_falseOut_valid,
      falseOut_ready => cond_br206_falseOut_ready
    );

  sink1 : entity work.sink_dataless(arch)
    port map(
      ins_valid => cond_br206_trueOut_valid,
      ins_ready => cond_br206_trueOut_ready,
      clk => clk,
      rst => rst
    );

  cond_br207 : entity work.cond_br(arch) generic map(32)
    port map(
      condition => fork51_outs_29,
      condition_valid => fork51_outs_29_valid,
      condition_ready => fork51_outs_29_ready,
      data => buffer37_outs,
      data_valid => buffer37_outs_valid,
      data_ready => buffer37_outs_ready,
      clk => clk,
      rst => rst,
      trueOut => cond_br207_trueOut,
      trueOut_valid => cond_br207_trueOut_valid,
      trueOut_ready => cond_br207_trueOut_ready,
      falseOut => cond_br207_falseOut,
      falseOut_valid => cond_br207_falseOut_valid,
      falseOut_ready => cond_br207_falseOut_ready
    );

  buffer37 : entity work.tfifo(arch) generic map(1, 32)
    port map(
      ins => fork10_outs_1,
      ins_valid => fork10_outs_1_valid,
      ins_ready => fork10_outs_1_ready,
      clk => clk,
      rst => rst,
      outs => buffer37_outs,
      outs_valid => buffer37_outs_valid,
      outs_ready => buffer37_outs_ready
    );

  sink2 : entity work.sink(arch) generic map(32)
    port map(
      ins => cond_br207_falseOut,
      ins_valid => cond_br207_falseOut_valid,
      ins_ready => cond_br207_falseOut_ready,
      clk => clk,
      rst => rst
    );

  cond_br208 : entity work.cond_br_dataless(arch)
    port map(
      condition => buffer38_outs,
      condition_valid => buffer38_outs_valid,
      condition_ready => buffer38_outs_ready,
      data_valid => fork45_outs_1_valid,
      data_ready => fork45_outs_1_ready,
      clk => clk,
      rst => rst,
      trueOut_valid => cond_br208_trueOut_valid,
      trueOut_ready => cond_br208_trueOut_ready,
      falseOut_valid => cond_br208_falseOut_valid,
      falseOut_ready => cond_br208_falseOut_ready
    );

  buffer38 : entity work.tfifo(arch) generic map(1, 1)
    port map(
      ins => fork51_outs_28,
      ins_valid => fork51_outs_28_valid,
      ins_ready => fork51_outs_28_ready,
      clk => clk,
      rst => rst,
      outs => buffer38_outs,
      outs_valid => buffer38_outs_valid,
      outs_ready => buffer38_outs_ready
    );

  sink3 : entity work.sink_dataless(arch)
    port map(
      ins_valid => cond_br208_trueOut_valid,
      ins_ready => cond_br208_trueOut_ready,
      clk => clk,
      rst => rst
    );

  cond_br209 : entity work.cond_br(arch) generic map(11)
    port map(
      condition => fork51_outs_1,
      condition_valid => fork51_outs_1_valid,
      condition_ready => fork51_outs_1_ready,
      data => fork7_outs_0,
      data_valid => fork7_outs_0_valid,
      data_ready => fork7_outs_0_ready,
      clk => clk,
      rst => rst,
      trueOut => cond_br209_trueOut,
      trueOut_valid => cond_br209_trueOut_valid,
      trueOut_ready => cond_br209_trueOut_ready,
      falseOut => cond_br209_falseOut,
      falseOut_valid => cond_br209_falseOut_valid,
      falseOut_ready => cond_br209_falseOut_ready
    );

  sink4 : entity work.sink(arch) generic map(11)
    port map(
      ins => cond_br209_falseOut,
      ins_valid => cond_br209_falseOut_valid,
      ins_ready => cond_br209_falseOut_ready,
      clk => clk,
      rst => rst
    );

  cond_br210 : entity work.cond_br_dataless(arch)
    port map(
      condition => fork51_outs_27,
      condition_valid => fork51_outs_27_valid,
      condition_ready => fork51_outs_27_ready,
      data_valid => fork38_outs_1_valid,
      data_ready => fork38_outs_1_ready,
      clk => clk,
      rst => rst,
      trueOut_valid => cond_br210_trueOut_valid,
      trueOut_ready => cond_br210_trueOut_ready,
      falseOut_valid => cond_br210_falseOut_valid,
      falseOut_ready => cond_br210_falseOut_ready
    );

  sink5 : entity work.sink_dataless(arch)
    port map(
      ins_valid => cond_br210_trueOut_valid,
      ins_ready => cond_br210_trueOut_ready,
      clk => clk,
      rst => rst
    );

  cond_br211 : entity work.cond_br(arch) generic map(32)
    port map(
      condition => fork51_outs_26,
      condition_valid => fork51_outs_26_valid,
      condition_ready => fork51_outs_26_ready,
      data => init89_outs,
      data_valid => init89_outs_valid,
      data_ready => init89_outs_ready,
      clk => clk,
      rst => rst,
      trueOut => cond_br211_trueOut,
      trueOut_valid => cond_br211_trueOut_valid,
      trueOut_ready => cond_br211_trueOut_ready,
      falseOut => cond_br211_falseOut,
      falseOut_valid => cond_br211_falseOut_valid,
      falseOut_ready => cond_br211_falseOut_ready
    );

  sink6 : entity work.sink(arch) generic map(32)
    port map(
      ins => cond_br211_trueOut,
      ins_valid => cond_br211_trueOut_valid,
      ins_ready => cond_br211_trueOut_ready,
      clk => clk,
      rst => rst
    );

  cond_br212 : entity work.cond_br(arch) generic map(8)
    port map(
      condition => fork51_outs_6,
      condition_valid => fork51_outs_6_valid,
      condition_ready => fork51_outs_6_ready,
      data => fork44_outs_0,
      data_valid => fork44_outs_0_valid,
      data_ready => fork44_outs_0_ready,
      clk => clk,
      rst => rst,
      trueOut => cond_br212_trueOut,
      trueOut_valid => cond_br212_trueOut_valid,
      trueOut_ready => cond_br212_trueOut_ready,
      falseOut => cond_br212_falseOut,
      falseOut_valid => cond_br212_falseOut_valid,
      falseOut_ready => cond_br212_falseOut_ready
    );

  sink7 : entity work.sink(arch) generic map(8)
    port map(
      ins => cond_br212_trueOut,
      ins_valid => cond_br212_trueOut_valid,
      ins_ready => cond_br212_trueOut_ready,
      clk => clk,
      rst => rst
    );

  cond_br213 : entity work.cond_br(arch) generic map(32)
    port map(
      condition => fork51_outs_25,
      condition_valid => fork51_outs_25_valid,
      condition_ready => fork51_outs_25_ready,
      data => fork6_outs_1,
      data_valid => fork6_outs_1_valid,
      data_ready => fork6_outs_1_ready,
      clk => clk,
      rst => rst,
      trueOut => cond_br213_trueOut,
      trueOut_valid => cond_br213_trueOut_valid,
      trueOut_ready => cond_br213_trueOut_ready,
      falseOut => cond_br213_falseOut,
      falseOut_valid => cond_br213_falseOut_valid,
      falseOut_ready => cond_br213_falseOut_ready
    );

  sink8 : entity work.sink(arch) generic map(32)
    port map(
      ins => cond_br213_falseOut,
      ins_valid => cond_br213_falseOut_valid,
      ins_ready => cond_br213_falseOut_ready,
      clk => clk,
      rst => rst
    );

  cond_br214 : entity work.cond_br_dataless(arch)
    port map(
      condition => fork51_outs_24,
      condition_valid => fork51_outs_24_valid,
      condition_ready => fork51_outs_24_ready,
      data_valid => init91_outs_valid,
      data_ready => init91_outs_ready,
      clk => clk,
      rst => rst,
      trueOut_valid => cond_br214_trueOut_valid,
      trueOut_ready => cond_br214_trueOut_ready,
      falseOut_valid => cond_br214_falseOut_valid,
      falseOut_ready => cond_br214_falseOut_ready
    );

  sink9 : entity work.sink_dataless(arch)
    port map(
      ins_valid => cond_br214_trueOut_valid,
      ins_ready => cond_br214_trueOut_ready,
      clk => clk,
      rst => rst
    );

  cond_br215 : entity work.cond_br_dataless(arch)
    port map(
      condition => fork51_outs_23,
      condition_valid => fork51_outs_23_valid,
      condition_ready => fork51_outs_23_ready,
      data_valid => fork21_outs_1_valid,
      data_ready => fork21_outs_1_ready,
      clk => clk,
      rst => rst,
      trueOut_valid => cond_br215_trueOut_valid,
      trueOut_ready => cond_br215_trueOut_ready,
      falseOut_valid => cond_br215_falseOut_valid,
      falseOut_ready => cond_br215_falseOut_ready
    );

  sink10 : entity work.sink_dataless(arch)
    port map(
      ins_valid => cond_br215_trueOut_valid,
      ins_ready => cond_br215_trueOut_ready,
      clk => clk,
      rst => rst
    );

  cond_br216 : entity work.cond_br_dataless(arch)
    port map(
      condition => fork51_outs_22,
      condition_valid => fork51_outs_22_valid,
      condition_ready => fork51_outs_22_ready,
      data_valid => fork22_outs_1_valid,
      data_ready => fork22_outs_1_ready,
      clk => clk,
      rst => rst,
      trueOut_valid => cond_br216_trueOut_valid,
      trueOut_ready => cond_br216_trueOut_ready,
      falseOut_valid => cond_br216_falseOut_valid,
      falseOut_ready => cond_br216_falseOut_ready
    );

  sink11 : entity work.sink_dataless(arch)
    port map(
      ins_valid => cond_br216_trueOut_valid,
      ins_ready => cond_br216_trueOut_ready,
      clk => clk,
      rst => rst
    );

  cond_br217 : entity work.cond_br(arch) generic map(32)
    port map(
      condition => fork51_outs_21,
      condition_valid => fork51_outs_21_valid,
      condition_ready => fork51_outs_21_ready,
      data => fork9_outs_1,
      data_valid => fork9_outs_1_valid,
      data_ready => fork9_outs_1_ready,
      clk => clk,
      rst => rst,
      trueOut => cond_br217_trueOut,
      trueOut_valid => cond_br217_trueOut_valid,
      trueOut_ready => cond_br217_trueOut_ready,
      falseOut => cond_br217_falseOut,
      falseOut_valid => cond_br217_falseOut_valid,
      falseOut_ready => cond_br217_falseOut_ready
    );

  sink12 : entity work.sink(arch) generic map(32)
    port map(
      ins => cond_br217_falseOut,
      ins_valid => cond_br217_falseOut_valid,
      ins_ready => cond_br217_falseOut_ready,
      clk => clk,
      rst => rst
    );

  cond_br218 : entity work.cond_br(arch) generic map(11)
    port map(
      condition => fork51_outs_3,
      condition_valid => fork51_outs_3_valid,
      condition_ready => fork51_outs_3_ready,
      data => fork13_outs_0,
      data_valid => fork13_outs_0_valid,
      data_ready => fork13_outs_0_ready,
      clk => clk,
      rst => rst,
      trueOut => cond_br218_trueOut,
      trueOut_valid => cond_br218_trueOut_valid,
      trueOut_ready => cond_br218_trueOut_ready,
      falseOut => cond_br218_falseOut,
      falseOut_valid => cond_br218_falseOut_valid,
      falseOut_ready => cond_br218_falseOut_ready
    );

  sink13 : entity work.sink(arch) generic map(11)
    port map(
      ins => cond_br218_falseOut,
      ins_valid => cond_br218_falseOut_valid,
      ins_ready => cond_br218_falseOut_ready,
      clk => clk,
      rst => rst
    );

  cond_br219 : entity work.cond_br_dataless(arch)
    port map(
      condition => fork51_outs_20,
      condition_valid => fork51_outs_20_valid,
      condition_ready => fork51_outs_20_ready,
      data_valid => init88_outs_valid,
      data_ready => init88_outs_ready,
      clk => clk,
      rst => rst,
      trueOut_valid => cond_br219_trueOut_valid,
      trueOut_ready => cond_br219_trueOut_ready,
      falseOut_valid => cond_br219_falseOut_valid,
      falseOut_ready => cond_br219_falseOut_ready
    );

  sink14 : entity work.sink_dataless(arch)
    port map(
      ins_valid => cond_br219_trueOut_valid,
      ins_ready => cond_br219_trueOut_ready,
      clk => clk,
      rst => rst
    );

  cond_br220 : entity work.cond_br(arch) generic map(9)
    port map(
      condition => fork51_outs_7,
      condition_valid => fork51_outs_7_valid,
      condition_ready => fork51_outs_7_ready,
      data => fork36_outs_0,
      data_valid => fork36_outs_0_valid,
      data_ready => fork36_outs_0_ready,
      clk => clk,
      rst => rst,
      trueOut => cond_br220_trueOut,
      trueOut_valid => cond_br220_trueOut_valid,
      trueOut_ready => cond_br220_trueOut_ready,
      falseOut => cond_br220_falseOut,
      falseOut_valid => cond_br220_falseOut_valid,
      falseOut_ready => cond_br220_falseOut_ready
    );

  sink15 : entity work.sink(arch) generic map(9)
    port map(
      ins => cond_br220_trueOut,
      ins_valid => cond_br220_trueOut_valid,
      ins_ready => cond_br220_trueOut_ready,
      clk => clk,
      rst => rst
    );

  cond_br221 : entity work.cond_br_dataless(arch)
    port map(
      condition => buffer57_outs,
      condition_valid => buffer57_outs_valid,
      condition_ready => buffer57_outs_ready,
      data_valid => fork37_outs_1_valid,
      data_ready => fork37_outs_1_ready,
      clk => clk,
      rst => rst,
      trueOut_valid => cond_br221_trueOut_valid,
      trueOut_ready => cond_br221_trueOut_ready,
      falseOut_valid => cond_br221_falseOut_valid,
      falseOut_ready => cond_br221_falseOut_ready
    );

  buffer57 : entity work.tfifo(arch) generic map(1, 1)
    port map(
      ins => fork51_outs_19,
      ins_valid => fork51_outs_19_valid,
      ins_ready => fork51_outs_19_ready,
      clk => clk,
      rst => rst,
      outs => buffer57_outs,
      outs_valid => buffer57_outs_valid,
      outs_ready => buffer57_outs_ready
    );

  sink16 : entity work.sink_dataless(arch)
    port map(
      ins_valid => cond_br221_trueOut_valid,
      ins_ready => cond_br221_trueOut_ready,
      clk => clk,
      rst => rst
    );

  cond_br222 : entity work.cond_br(arch) generic map(11)
    port map(
      condition => fork51_outs_2,
      condition_valid => fork51_outs_2_valid,
      condition_ready => fork51_outs_2_ready,
      data => fork8_outs_0,
      data_valid => fork8_outs_0_valid,
      data_ready => fork8_outs_0_ready,
      clk => clk,
      rst => rst,
      trueOut => cond_br222_trueOut,
      trueOut_valid => cond_br222_trueOut_valid,
      trueOut_ready => cond_br222_trueOut_ready,
      falseOut => cond_br222_falseOut,
      falseOut_valid => cond_br222_falseOut_valid,
      falseOut_ready => cond_br222_falseOut_ready
    );

  sink17 : entity work.sink(arch) generic map(11)
    port map(
      ins => cond_br222_falseOut,
      ins_valid => cond_br222_falseOut_valid,
      ins_ready => cond_br222_falseOut_ready,
      clk => clk,
      rst => rst
    );

  cond_br223 : entity work.cond_br_dataless(arch)
    port map(
      condition => fork51_outs_18,
      condition_valid => fork51_outs_18_valid,
      condition_ready => fork51_outs_18_ready,
      data_valid => init85_outs_valid,
      data_ready => init85_outs_ready,
      clk => clk,
      rst => rst,
      trueOut_valid => cond_br223_trueOut_valid,
      trueOut_ready => cond_br223_trueOut_ready,
      falseOut_valid => cond_br223_falseOut_valid,
      falseOut_ready => cond_br223_falseOut_ready
    );

  sink18 : entity work.sink_dataless(arch)
    port map(
      ins_valid => cond_br223_trueOut_valid,
      ins_ready => cond_br223_trueOut_ready,
      clk => clk,
      rst => rst
    );

  cond_br224 : entity work.cond_br(arch) generic map(32)
    port map(
      condition => fork51_outs_17,
      condition_valid => fork51_outs_17_valid,
      condition_ready => fork51_outs_17_ready,
      data => init80_outs,
      data_valid => init80_outs_valid,
      data_ready => init80_outs_ready,
      clk => clk,
      rst => rst,
      trueOut => cond_br224_trueOut,
      trueOut_valid => cond_br224_trueOut_valid,
      trueOut_ready => cond_br224_trueOut_ready,
      falseOut => cond_br224_falseOut,
      falseOut_valid => cond_br224_falseOut_valid,
      falseOut_ready => cond_br224_falseOut_ready
    );

  sink19 : entity work.sink(arch) generic map(32)
    port map(
      ins => cond_br224_trueOut,
      ins_valid => cond_br224_trueOut_valid,
      ins_ready => cond_br224_trueOut_ready,
      clk => clk,
      rst => rst
    );

  cond_br225 : entity work.cond_br(arch) generic map(32)
    port map(
      condition => fork51_outs_16,
      condition_valid => fork51_outs_16_valid,
      condition_ready => fork51_outs_16_ready,
      data => init83_outs,
      data_valid => init83_outs_valid,
      data_ready => init83_outs_ready,
      clk => clk,
      rst => rst,
      trueOut => cond_br225_trueOut,
      trueOut_valid => cond_br225_trueOut_valid,
      trueOut_ready => cond_br225_trueOut_ready,
      falseOut => cond_br225_falseOut,
      falseOut_valid => cond_br225_falseOut_valid,
      falseOut_ready => cond_br225_falseOut_ready
    );

  sink20 : entity work.sink(arch) generic map(32)
    port map(
      ins => cond_br225_trueOut,
      ins_valid => cond_br225_trueOut_valid,
      ins_ready => cond_br225_trueOut_ready,
      clk => clk,
      rst => rst
    );

  cond_br226 : entity work.cond_br_dataless(arch)
    port map(
      condition => fork51_outs_15,
      condition_valid => fork51_outs_15_valid,
      condition_ready => fork51_outs_15_ready,
      data_valid => fork28_outs_1_valid,
      data_ready => fork28_outs_1_ready,
      clk => clk,
      rst => rst,
      trueOut_valid => cond_br226_trueOut_valid,
      trueOut_ready => cond_br226_trueOut_ready,
      falseOut_valid => cond_br226_falseOut_valid,
      falseOut_ready => cond_br226_falseOut_ready
    );

  sink21 : entity work.sink_dataless(arch)
    port map(
      ins_valid => cond_br226_trueOut_valid,
      ins_ready => cond_br226_trueOut_ready,
      clk => clk,
      rst => rst
    );

  cond_br227 : entity work.cond_br(arch) generic map(32)
    port map(
      condition => fork51_outs_14,
      condition_valid => fork51_outs_14_valid,
      condition_ready => fork51_outs_14_ready,
      data => init86_outs,
      data_valid => init86_outs_valid,
      data_ready => init86_outs_ready,
      clk => clk,
      rst => rst,
      trueOut => cond_br227_trueOut,
      trueOut_valid => cond_br227_trueOut_valid,
      trueOut_ready => cond_br227_trueOut_ready,
      falseOut => cond_br227_falseOut,
      falseOut_valid => cond_br227_falseOut_valid,
      falseOut_ready => cond_br227_falseOut_ready
    );

  sink22 : entity work.sink(arch) generic map(32)
    port map(
      ins => cond_br227_trueOut,
      ins_valid => cond_br227_trueOut_valid,
      ins_ready => cond_br227_trueOut_ready,
      clk => clk,
      rst => rst
    );

  cond_br228 : entity work.cond_br_dataless(arch)
    port map(
      condition => fork51_outs_13,
      condition_valid => fork51_outs_13_valid,
      condition_ready => fork51_outs_13_ready,
      data_valid => fork5_outs_12_valid,
      data_ready => fork5_outs_12_ready,
      clk => clk,
      rst => rst,
      trueOut_valid => cond_br228_trueOut_valid,
      trueOut_ready => cond_br228_trueOut_ready,
      falseOut_valid => cond_br228_falseOut_valid,
      falseOut_ready => cond_br228_falseOut_ready
    );

  sink23 : entity work.sink_dataless(arch)
    port map(
      ins_valid => cond_br228_falseOut_valid,
      ins_ready => cond_br228_falseOut_ready,
      clk => clk,
      rst => rst
    );

  cond_br229 : entity work.cond_br_dataless(arch)
    port map(
      condition => buffer66_outs,
      condition_valid => buffer66_outs_valid,
      condition_ready => buffer66_outs_ready,
      data_valid => fork46_outs_1_valid,
      data_ready => fork46_outs_1_ready,
      clk => clk,
      rst => rst,
      trueOut_valid => cond_br229_trueOut_valid,
      trueOut_ready => cond_br229_trueOut_ready,
      falseOut_valid => cond_br229_falseOut_valid,
      falseOut_ready => cond_br229_falseOut_ready
    );

  buffer66 : entity work.tfifo(arch) generic map(1, 1)
    port map(
      ins => fork51_outs_12,
      ins_valid => fork51_outs_12_valid,
      ins_ready => fork51_outs_12_ready,
      clk => clk,
      rst => rst,
      outs => buffer66_outs,
      outs_valid => buffer66_outs_valid,
      outs_ready => buffer66_outs_ready
    );

  sink24 : entity work.sink_dataless(arch)
    port map(
      ins_valid => cond_br229_trueOut_valid,
      ins_ready => cond_br229_trueOut_ready,
      clk => clk,
      rst => rst
    );

  cond_br230 : entity work.cond_br(arch) generic map(8)
    port map(
      condition => fork51_outs_8,
      condition_valid => fork51_outs_8_valid,
      condition_ready => fork51_outs_8_ready,
      data => buffer68_outs,
      data_valid => buffer68_outs_valid,
      data_ready => buffer68_outs_ready,
      clk => clk,
      rst => rst,
      trueOut => cond_br230_trueOut,
      trueOut_valid => cond_br230_trueOut_valid,
      trueOut_ready => cond_br230_trueOut_ready,
      falseOut => cond_br230_falseOut,
      falseOut_valid => cond_br230_falseOut_valid,
      falseOut_ready => cond_br230_falseOut_ready
    );

  buffer68 : entity work.tfifo(arch) generic map(1, 8)
    port map(
      ins => fork27_outs_0,
      ins_valid => fork27_outs_0_valid,
      ins_ready => fork27_outs_0_ready,
      clk => clk,
      rst => rst,
      outs => buffer68_outs,
      outs_valid => buffer68_outs_valid,
      outs_ready => buffer68_outs_ready
    );

  sink25 : entity work.sink(arch) generic map(8)
    port map(
      ins => cond_br230_trueOut,
      ins_valid => cond_br230_trueOut_valid,
      ins_ready => cond_br230_trueOut_ready,
      clk => clk,
      rst => rst
    );

  cond_br231 : entity work.cond_br_dataless(arch)
    port map(
      condition => fork51_outs_11,
      condition_valid => fork51_outs_11_valid,
      condition_ready => fork51_outs_11_ready,
      data_valid => init82_outs_valid,
      data_ready => init82_outs_ready,
      clk => clk,
      rst => rst,
      trueOut_valid => cond_br231_trueOut_valid,
      trueOut_ready => cond_br231_trueOut_ready,
      falseOut_valid => cond_br231_falseOut_valid,
      falseOut_ready => cond_br231_falseOut_ready
    );

  sink26 : entity work.sink_dataless(arch)
    port map(
      ins_valid => cond_br231_trueOut_valid,
      ins_ready => cond_br231_trueOut_ready,
      clk => clk,
      rst => rst
    );

  cond_br232 : entity work.cond_br(arch) generic map(32)
    port map(
      condition => fork51_outs_10,
      condition_valid => fork51_outs_10_valid,
      condition_ready => fork51_outs_10_ready,
      data => fork20_outs_1,
      data_valid => fork20_outs_1_valid,
      data_ready => fork20_outs_1_ready,
      clk => clk,
      rst => rst,
      trueOut => cond_br232_trueOut,
      trueOut_valid => cond_br232_trueOut_valid,
      trueOut_ready => cond_br232_trueOut_ready,
      falseOut => cond_br232_falseOut,
      falseOut_valid => cond_br232_falseOut_valid,
      falseOut_ready => cond_br232_falseOut_ready
    );

  sink27 : entity work.sink(arch) generic map(32)
    port map(
      ins => cond_br232_trueOut,
      ins_valid => cond_br232_trueOut_valid,
      ins_ready => cond_br232_trueOut_ready,
      clk => clk,
      rst => rst
    );

  cond_br233 : entity work.cond_br(arch) generic map(11)
    port map(
      condition => fork51_outs_4,
      condition_valid => fork51_outs_4_valid,
      condition_ready => fork51_outs_4_ready,
      data => fork12_outs_0,
      data_valid => fork12_outs_0_valid,
      data_ready => fork12_outs_0_ready,
      clk => clk,
      rst => rst,
      trueOut => cond_br233_trueOut,
      trueOut_valid => cond_br233_trueOut_valid,
      trueOut_ready => cond_br233_trueOut_ready,
      falseOut => cond_br233_falseOut,
      falseOut_valid => cond_br233_falseOut_valid,
      falseOut_ready => cond_br233_falseOut_ready
    );

  sink28 : entity work.sink(arch) generic map(11)
    port map(
      ins => cond_br233_falseOut,
      ins_valid => cond_br233_falseOut_valid,
      ins_ready => cond_br233_falseOut_ready,
      clk => clk,
      rst => rst
    );

  init40 : entity work.tehb_init(arch) generic map(1, 0)
    port map(
      ins => fork51_outs_9,
      ins_valid => fork51_outs_9_valid,
      ins_ready => fork51_outs_9_ready,
      clk => clk,
      rst => rst,
      outs => init40_outs,
      outs_valid => init40_outs_valid,
      outs_ready => init40_outs_ready
    );

  fork4 : entity work.handshake_fork(arch) generic map(9, 1)
    port map(
      ins => init40_outs,
      ins_valid => init40_outs_valid,
      ins_ready => init40_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork4_outs_0,
      outs(1) => fork4_outs_1,
      outs(2) => fork4_outs_2,
      outs(3) => fork4_outs_3,
      outs(4) => fork4_outs_4,
      outs(5) => fork4_outs_5,
      outs(6) => fork4_outs_6,
      outs(7) => fork4_outs_7,
      outs(8) => fork4_outs_8,
      outs_valid(0) => fork4_outs_0_valid,
      outs_valid(1) => fork4_outs_1_valid,
      outs_valid(2) => fork4_outs_2_valid,
      outs_valid(3) => fork4_outs_3_valid,
      outs_valid(4) => fork4_outs_4_valid,
      outs_valid(5) => fork4_outs_5_valid,
      outs_valid(6) => fork4_outs_6_valid,
      outs_valid(7) => fork4_outs_7_valid,
      outs_valid(8) => fork4_outs_8_valid,
      outs_ready(0) => fork4_outs_0_ready,
      outs_ready(1) => fork4_outs_1_ready,
      outs_ready(2) => fork4_outs_2_ready,
      outs_ready(3) => fork4_outs_3_ready,
      outs_ready(4) => fork4_outs_4_ready,
      outs_ready(5) => fork4_outs_5_ready,
      outs_ready(6) => fork4_outs_6_ready,
      outs_ready(7) => fork4_outs_7_ready,
      outs_ready(8) => fork4_outs_8_ready
    );

  buffer12 : entity work.tehb_dataless(arch)
    port map(
      ins_valid => mux37_outs_valid,
      ins_ready => mux37_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer12_outs_valid,
      outs_ready => buffer12_outs_ready
    );

  mux45 : entity work.mux_dataless(arch) generic map(2, 1)
    port map(
      index => fork4_outs_8,
      index_valid => fork4_outs_8_valid,
      index_ready => fork4_outs_8_ready,
      ins_valid(0) => buffer12_outs_valid,
      ins_valid(1) => cond_br228_trueOut_valid,
      ins_ready(0) => buffer12_outs_ready,
      ins_ready(1) => cond_br228_trueOut_ready,
      clk => clk,
      rst => rst,
      outs_valid => mux45_outs_valid,
      outs_ready => mux45_outs_ready
    );

  buffer14 : entity work.oehb_dataless(arch)
    port map(
      ins_valid => mux45_outs_valid,
      ins_ready => mux45_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer14_outs_valid,
      outs_ready => buffer14_outs_ready
    );

  buffer15 : entity work.tehb_dataless(arch)
    port map(
      ins_valid => buffer14_outs_valid,
      ins_ready => buffer14_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer15_outs_valid,
      outs_ready => buffer15_outs_ready
    );

  fork5 : entity work.fork_dataless(arch) generic map(13)
    port map(
      ins_valid => buffer15_outs_valid,
      ins_ready => buffer15_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid(0) => fork5_outs_0_valid,
      outs_valid(1) => fork5_outs_1_valid,
      outs_valid(2) => fork5_outs_2_valid,
      outs_valid(3) => fork5_outs_3_valid,
      outs_valid(4) => fork5_outs_4_valid,
      outs_valid(5) => fork5_outs_5_valid,
      outs_valid(6) => fork5_outs_6_valid,
      outs_valid(7) => fork5_outs_7_valid,
      outs_valid(8) => fork5_outs_8_valid,
      outs_valid(9) => fork5_outs_9_valid,
      outs_valid(10) => fork5_outs_10_valid,
      outs_valid(11) => fork5_outs_11_valid,
      outs_valid(12) => fork5_outs_12_valid,
      outs_ready(0) => fork5_outs_0_ready,
      outs_ready(1) => fork5_outs_1_ready,
      outs_ready(2) => fork5_outs_2_ready,
      outs_ready(3) => fork5_outs_3_ready,
      outs_ready(4) => fork5_outs_4_ready,
      outs_ready(5) => fork5_outs_5_ready,
      outs_ready(6) => fork5_outs_6_ready,
      outs_ready(7) => fork5_outs_7_ready,
      outs_ready(8) => fork5_outs_8_ready,
      outs_ready(9) => fork5_outs_9_ready,
      outs_ready(10) => fork5_outs_10_ready,
      outs_ready(11) => fork5_outs_11_ready,
      outs_ready(12) => fork5_outs_12_ready
    );

  mux48 : entity work.mux(arch) generic map(2, 32, 1)
    port map(
      index => fork4_outs_7,
      index_valid => fork4_outs_7_valid,
      index_ready => fork4_outs_7_ready,
      ins(0) => mux21_outs,
      ins(1) => cond_br213_trueOut,
      ins_valid(0) => mux21_outs_valid,
      ins_valid(1) => cond_br213_trueOut_valid,
      ins_ready(0) => mux21_outs_ready,
      ins_ready(1) => cond_br213_trueOut_ready,
      clk => clk,
      rst => rst,
      outs => mux48_outs,
      outs_valid => mux48_outs_valid,
      outs_ready => mux48_outs_ready
    );

  buffer16 : entity work.oehb(arch) generic map(32)
    port map(
      ins => mux48_outs,
      ins_valid => mux48_outs_valid,
      ins_ready => mux48_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer16_outs,
      outs_valid => buffer16_outs_valid,
      outs_ready => buffer16_outs_ready
    );

  buffer17 : entity work.tehb(arch) generic map(32)
    port map(
      ins => buffer16_outs,
      ins_valid => buffer16_outs_valid,
      ins_ready => buffer16_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer17_outs,
      outs_valid => buffer17_outs_valid,
      outs_ready => buffer17_outs_ready
    );

  fork6 : entity work.handshake_fork(arch) generic map(2, 32)
    port map(
      ins => buffer17_outs,
      ins_valid => buffer17_outs_valid,
      ins_ready => buffer17_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork6_outs_0,
      outs(1) => fork6_outs_1,
      outs_valid(0) => fork6_outs_0_valid,
      outs_valid(1) => fork6_outs_1_valid,
      outs_ready(0) => fork6_outs_0_ready,
      outs_ready(1) => fork6_outs_1_ready
    );

  mux51 : entity work.mux(arch) generic map(2, 11, 1)
    port map(
      index => fork4_outs_0,
      index_valid => fork4_outs_0_valid,
      index_ready => fork4_outs_0_ready,
      ins(0) => mux9_outs,
      ins(1) => cond_br209_trueOut,
      ins_valid(0) => mux9_outs_valid,
      ins_valid(1) => cond_br209_trueOut_valid,
      ins_ready(0) => mux9_outs_ready,
      ins_ready(1) => cond_br209_trueOut_ready,
      clk => clk,
      rst => rst,
      outs => mux51_outs,
      outs_valid => mux51_outs_valid,
      outs_ready => mux51_outs_ready
    );

  buffer18 : entity work.oehb(arch) generic map(11)
    port map(
      ins => mux51_outs,
      ins_valid => mux51_outs_valid,
      ins_ready => mux51_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer18_outs,
      outs_valid => buffer18_outs_valid,
      outs_ready => buffer18_outs_ready
    );

  buffer19 : entity work.tehb(arch) generic map(11)
    port map(
      ins => buffer18_outs,
      ins_valid => buffer18_outs_valid,
      ins_ready => buffer18_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer19_outs,
      outs_valid => buffer19_outs_valid,
      outs_ready => buffer19_outs_ready
    );

  fork7 : entity work.handshake_fork(arch) generic map(2, 11)
    port map(
      ins => buffer19_outs,
      ins_valid => buffer19_outs_valid,
      ins_ready => buffer19_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork7_outs_0,
      outs(1) => fork7_outs_1,
      outs_valid(0) => fork7_outs_0_valid,
      outs_valid(1) => fork7_outs_1_valid,
      outs_ready(0) => fork7_outs_0_ready,
      outs_ready(1) => fork7_outs_1_ready
    );

  extsi22 : entity work.extsi(arch) generic map(11, 32)
    port map(
      ins => fork7_outs_1,
      ins_valid => fork7_outs_1_valid,
      ins_ready => fork7_outs_1_ready,
      clk => clk,
      rst => rst,
      outs => extsi22_outs,
      outs_valid => extsi22_outs_valid,
      outs_ready => extsi22_outs_ready
    );

  mux52 : entity work.mux(arch) generic map(2, 11, 1)
    port map(
      index => fork4_outs_1,
      index_valid => fork4_outs_1_valid,
      index_ready => fork4_outs_1_ready,
      ins(0) => mux10_outs,
      ins(1) => cond_br222_trueOut,
      ins_valid(0) => mux10_outs_valid,
      ins_valid(1) => cond_br222_trueOut_valid,
      ins_ready(0) => mux10_outs_ready,
      ins_ready(1) => cond_br222_trueOut_ready,
      clk => clk,
      rst => rst,
      outs => mux52_outs,
      outs_valid => mux52_outs_valid,
      outs_ready => mux52_outs_ready
    );

  buffer20 : entity work.oehb(arch) generic map(11)
    port map(
      ins => mux52_outs,
      ins_valid => mux52_outs_valid,
      ins_ready => mux52_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer20_outs,
      outs_valid => buffer20_outs_valid,
      outs_ready => buffer20_outs_ready
    );

  buffer21 : entity work.tehb(arch) generic map(11)
    port map(
      ins => buffer20_outs,
      ins_valid => buffer20_outs_valid,
      ins_ready => buffer20_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer21_outs,
      outs_valid => buffer21_outs_valid,
      outs_ready => buffer21_outs_ready
    );

  fork8 : entity work.handshake_fork(arch) generic map(2, 11)
    port map(
      ins => buffer21_outs,
      ins_valid => buffer21_outs_valid,
      ins_ready => buffer21_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork8_outs_0,
      outs(1) => fork8_outs_1,
      outs_valid(0) => fork8_outs_0_valid,
      outs_valid(1) => fork8_outs_1_valid,
      outs_ready(0) => fork8_outs_0_ready,
      outs_ready(1) => fork8_outs_1_ready
    );

  extsi23 : entity work.extsi(arch) generic map(11, 32)
    port map(
      ins => fork8_outs_1,
      ins_valid => fork8_outs_1_valid,
      ins_ready => fork8_outs_1_ready,
      clk => clk,
      rst => rst,
      outs => extsi23_outs,
      outs_valid => extsi23_outs_valid,
      outs_ready => extsi23_outs_ready
    );

  mux54 : entity work.mux(arch) generic map(2, 32, 1)
    port map(
      index => fork4_outs_6,
      index_valid => fork4_outs_6_valid,
      index_ready => fork4_outs_6_ready,
      ins(0) => mux6_outs,
      ins(1) => cond_br217_trueOut,
      ins_valid(0) => mux6_outs_valid,
      ins_valid(1) => cond_br217_trueOut_valid,
      ins_ready(0) => mux6_outs_ready,
      ins_ready(1) => cond_br217_trueOut_ready,
      clk => clk,
      rst => rst,
      outs => mux54_outs,
      outs_valid => mux54_outs_valid,
      outs_ready => mux54_outs_ready
    );

  buffer22 : entity work.oehb(arch) generic map(32)
    port map(
      ins => mux54_outs,
      ins_valid => mux54_outs_valid,
      ins_ready => mux54_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer22_outs,
      outs_valid => buffer22_outs_valid,
      outs_ready => buffer22_outs_ready
    );

  buffer23 : entity work.tehb(arch) generic map(32)
    port map(
      ins => buffer22_outs,
      ins_valid => buffer22_outs_valid,
      ins_ready => buffer22_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer23_outs,
      outs_valid => buffer23_outs_valid,
      outs_ready => buffer23_outs_ready
    );

  fork9 : entity work.handshake_fork(arch) generic map(2, 32)
    port map(
      ins => buffer23_outs,
      ins_valid => buffer23_outs_valid,
      ins_ready => buffer23_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork9_outs_0,
      outs(1) => fork9_outs_1,
      outs_valid(0) => fork9_outs_0_valid,
      outs_valid(1) => fork9_outs_1_valid,
      outs_ready(0) => fork9_outs_0_ready,
      outs_ready(1) => fork9_outs_1_ready
    );

  mux56 : entity work.mux(arch) generic map(2, 32, 1)
    port map(
      index => fork4_outs_5,
      index_valid => fork4_outs_5_valid,
      index_ready => fork4_outs_5_ready,
      ins(0) => mux7_outs,
      ins(1) => cond_br207_trueOut,
      ins_valid(0) => mux7_outs_valid,
      ins_valid(1) => cond_br207_trueOut_valid,
      ins_ready(0) => mux7_outs_ready,
      ins_ready(1) => cond_br207_trueOut_ready,
      clk => clk,
      rst => rst,
      outs => mux56_outs,
      outs_valid => mux56_outs_valid,
      outs_ready => mux56_outs_ready
    );

  buffer24 : entity work.oehb(arch) generic map(32)
    port map(
      ins => mux56_outs,
      ins_valid => mux56_outs_valid,
      ins_ready => mux56_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer24_outs,
      outs_valid => buffer24_outs_valid,
      outs_ready => buffer24_outs_ready
    );

  buffer25 : entity work.tehb(arch) generic map(32)
    port map(
      ins => buffer24_outs,
      ins_valid => buffer24_outs_valid,
      ins_ready => buffer24_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer25_outs,
      outs_valid => buffer25_outs_valid,
      outs_ready => buffer25_outs_ready
    );

  fork10 : entity work.handshake_fork(arch) generic map(2, 32)
    port map(
      ins => buffer25_outs,
      ins_valid => buffer25_outs_valid,
      ins_ready => buffer25_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork10_outs_0,
      outs(1) => fork10_outs_1,
      outs_valid(0) => fork10_outs_0_valid,
      outs_valid(1) => fork10_outs_1_valid,
      outs_ready(0) => fork10_outs_0_ready,
      outs_ready(1) => fork10_outs_1_ready
    );

  mux57 : entity work.mux(arch) generic map(2, 32, 1)
    port map(
      index => fork4_outs_4,
      index_valid => fork4_outs_4_valid,
      index_ready => fork4_outs_4_ready,
      ins(0) => mux23_outs,
      ins(1) => cond_br205_trueOut,
      ins_valid(0) => mux23_outs_valid,
      ins_valid(1) => cond_br205_trueOut_valid,
      ins_ready(0) => mux23_outs_ready,
      ins_ready(1) => cond_br205_trueOut_ready,
      clk => clk,
      rst => rst,
      outs => mux57_outs,
      outs_valid => mux57_outs_valid,
      outs_ready => mux57_outs_ready
    );

  buffer26 : entity work.oehb(arch) generic map(32)
    port map(
      ins => mux57_outs,
      ins_valid => mux57_outs_valid,
      ins_ready => mux57_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer26_outs,
      outs_valid => buffer26_outs_valid,
      outs_ready => buffer26_outs_ready
    );

  buffer27 : entity work.tehb(arch) generic map(32)
    port map(
      ins => buffer26_outs,
      ins_valid => buffer26_outs_valid,
      ins_ready => buffer26_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer27_outs,
      outs_valid => buffer27_outs_valid,
      outs_ready => buffer27_outs_ready
    );

  fork11 : entity work.handshake_fork(arch) generic map(2, 32)
    port map(
      ins => buffer27_outs,
      ins_valid => buffer27_outs_valid,
      ins_ready => buffer27_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork11_outs_0,
      outs(1) => fork11_outs_1,
      outs_valid(0) => fork11_outs_0_valid,
      outs_valid(1) => fork11_outs_1_valid,
      outs_ready(0) => fork11_outs_0_ready,
      outs_ready(1) => fork11_outs_1_ready
    );

  mux58 : entity work.mux(arch) generic map(2, 11, 1)
    port map(
      index => fork4_outs_3,
      index_valid => fork4_outs_3_valid,
      index_ready => fork4_outs_3_ready,
      ins(0) => mux28_outs,
      ins(1) => cond_br233_trueOut,
      ins_valid(0) => mux28_outs_valid,
      ins_valid(1) => cond_br233_trueOut_valid,
      ins_ready(0) => mux28_outs_ready,
      ins_ready(1) => cond_br233_trueOut_ready,
      clk => clk,
      rst => rst,
      outs => mux58_outs,
      outs_valid => mux58_outs_valid,
      outs_ready => mux58_outs_ready
    );

  buffer28 : entity work.oehb(arch) generic map(11)
    port map(
      ins => mux58_outs,
      ins_valid => mux58_outs_valid,
      ins_ready => mux58_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer28_outs,
      outs_valid => buffer28_outs_valid,
      outs_ready => buffer28_outs_ready
    );

  buffer29 : entity work.tehb(arch) generic map(11)
    port map(
      ins => buffer28_outs,
      ins_valid => buffer28_outs_valid,
      ins_ready => buffer28_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer29_outs,
      outs_valid => buffer29_outs_valid,
      outs_ready => buffer29_outs_ready
    );

  fork12 : entity work.handshake_fork(arch) generic map(2, 11)
    port map(
      ins => buffer29_outs,
      ins_valid => buffer29_outs_valid,
      ins_ready => buffer29_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork12_outs_0,
      outs(1) => fork12_outs_1,
      outs_valid(0) => fork12_outs_0_valid,
      outs_valid(1) => fork12_outs_1_valid,
      outs_ready(0) => fork12_outs_0_ready,
      outs_ready(1) => fork12_outs_1_ready
    );

  extsi24 : entity work.extsi(arch) generic map(11, 32)
    port map(
      ins => fork12_outs_1,
      ins_valid => fork12_outs_1_valid,
      ins_ready => fork12_outs_1_ready,
      clk => clk,
      rst => rst,
      outs => extsi24_outs,
      outs_valid => extsi24_outs_valid,
      outs_ready => extsi24_outs_ready
    );

  mux60 : entity work.mux(arch) generic map(2, 11, 1)
    port map(
      index => fork4_outs_2,
      index_valid => fork4_outs_2_valid,
      index_ready => fork4_outs_2_ready,
      ins(0) => mux19_outs,
      ins(1) => cond_br218_trueOut,
      ins_valid(0) => mux19_outs_valid,
      ins_valid(1) => cond_br218_trueOut_valid,
      ins_ready(0) => mux19_outs_ready,
      ins_ready(1) => cond_br218_trueOut_ready,
      clk => clk,
      rst => rst,
      outs => mux60_outs,
      outs_valid => mux60_outs_valid,
      outs_ready => mux60_outs_ready
    );

  buffer30 : entity work.oehb(arch) generic map(11)
    port map(
      ins => mux60_outs,
      ins_valid => mux60_outs_valid,
      ins_ready => mux60_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer30_outs,
      outs_valid => buffer30_outs_valid,
      outs_ready => buffer30_outs_ready
    );

  buffer31 : entity work.tehb(arch) generic map(11)
    port map(
      ins => buffer30_outs,
      ins_valid => buffer30_outs_valid,
      ins_ready => buffer30_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer31_outs,
      outs_valid => buffer31_outs_valid,
      outs_ready => buffer31_outs_ready
    );

  fork13 : entity work.handshake_fork(arch) generic map(2, 11)
    port map(
      ins => buffer31_outs,
      ins_valid => buffer31_outs_valid,
      ins_ready => buffer31_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork13_outs_0,
      outs(1) => fork13_outs_1,
      outs_valid(0) => fork13_outs_0_valid,
      outs_valid(1) => fork13_outs_1_valid,
      outs_ready(0) => fork13_outs_0_ready,
      outs_ready(1) => fork13_outs_1_ready
    );

  extsi25 : entity work.extsi(arch) generic map(11, 32)
    port map(
      ins => fork13_outs_1,
      ins_valid => fork13_outs_1_valid,
      ins_ready => fork13_outs_1_ready,
      clk => clk,
      rst => rst,
      outs => extsi25_outs,
      outs_valid => extsi25_outs_valid,
      outs_ready => extsi25_outs_ready
    );

  unbundle3 : entity work.unbundle(arch) generic map(32)
    port map(
      ins => fork33_outs_0,
      ins_valid => fork33_outs_0_valid,
      ins_ready => fork33_outs_0_ready,
      clk => clk,
      rst => rst,
      outs_valid => unbundle3_outs_0_valid,
      outs_ready => unbundle3_outs_0_ready,
      outs => unbundle3_outs_1
    );

  unbundle4 : entity work.unbundle(arch) generic map(32)
    port map(
      ins => fork26_outs_0,
      ins_valid => fork26_outs_0_valid,
      ins_ready => fork26_outs_0_ready,
      clk => clk,
      rst => rst,
      outs_valid => unbundle4_outs_0_valid,
      outs_ready => unbundle4_outs_0_ready,
      outs => unbundle4_outs_1
    );

  unbundle5 : entity work.unbundle(arch) generic map(32)
    port map(
      ins => fork42_outs_0,
      ins_valid => fork42_outs_0_valid,
      ins_ready => fork42_outs_0_ready,
      clk => clk,
      rst => rst,
      outs_valid => unbundle5_outs_0_valid,
      outs_ready => unbundle5_outs_0_ready,
      outs => unbundle5_outs_1
    );

  mux1 : entity work.mux(arch) generic map(2, 8, 1)
    port map(
      index => fork16_outs_1,
      index_valid => fork16_outs_1_valid,
      index_ready => fork16_outs_1_ready,
      ins(0) => extsi20_outs,
      ins(1) => cond_br3_trueOut,
      ins_valid(0) => extsi20_outs_valid,
      ins_valid(1) => cond_br3_trueOut_valid,
      ins_ready(0) => extsi20_outs_ready,
      ins_ready(1) => cond_br3_trueOut_ready,
      clk => clk,
      rst => rst,
      outs => mux1_outs,
      outs_valid => mux1_outs_valid,
      outs_ready => mux1_outs_ready
    );

  buffer32 : entity work.oehb(arch) generic map(8)
    port map(
      ins => mux1_outs,
      ins_valid => mux1_outs_valid,
      ins_ready => mux1_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer32_outs,
      outs_valid => buffer32_outs_valid,
      outs_ready => buffer32_outs_ready
    );

  buffer33 : entity work.tehb(arch) generic map(8)
    port map(
      ins => buffer32_outs,
      ins_valid => buffer32_outs_valid,
      ins_ready => buffer32_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer33_outs,
      outs_valid => buffer33_outs_valid,
      outs_ready => buffer33_outs_ready
    );

  fork14 : entity work.handshake_fork(arch) generic map(5, 8)
    port map(
      ins => buffer33_outs,
      ins_valid => buffer33_outs_valid,
      ins_ready => buffer33_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork14_outs_0,
      outs(1) => fork14_outs_1,
      outs(2) => fork14_outs_2,
      outs(3) => fork14_outs_3,
      outs(4) => fork14_outs_4,
      outs_valid(0) => fork14_outs_0_valid,
      outs_valid(1) => fork14_outs_1_valid,
      outs_valid(2) => fork14_outs_2_valid,
      outs_valid(3) => fork14_outs_3_valid,
      outs_valid(4) => fork14_outs_4_valid,
      outs_ready(0) => fork14_outs_0_ready,
      outs_ready(1) => fork14_outs_1_ready,
      outs_ready(2) => fork14_outs_2_ready,
      outs_ready(3) => fork14_outs_3_ready,
      outs_ready(4) => fork14_outs_4_ready
    );

  extsi26 : entity work.extsi(arch) generic map(8, 9)
    port map(
      ins => fork14_outs_0,
      ins_valid => fork14_outs_0_valid,
      ins_ready => fork14_outs_0_ready,
      clk => clk,
      rst => rst,
      outs => extsi26_outs,
      outs_valid => extsi26_outs_valid,
      outs_ready => extsi26_outs_ready
    );

  extsi27 : entity work.extsi(arch) generic map(8, 9)
    port map(
      ins => fork14_outs_2,
      ins_valid => fork14_outs_2_valid,
      ins_ready => fork14_outs_2_ready,
      clk => clk,
      rst => rst,
      outs => extsi27_outs,
      outs_valid => extsi27_outs_valid,
      outs_ready => extsi27_outs_ready
    );

  extsi28 : entity work.extsi(arch) generic map(8, 32)
    port map(
      ins => fork14_outs_4,
      ins_valid => fork14_outs_4_valid,
      ins_ready => fork14_outs_4_ready,
      clk => clk,
      rst => rst,
      outs => extsi28_outs,
      outs_valid => extsi28_outs_valid,
      outs_ready => extsi28_outs_ready
    );

  fork15 : entity work.handshake_fork(arch) generic map(5, 32)
    port map(
      ins => extsi28_outs,
      ins_valid => extsi28_outs_valid,
      ins_ready => extsi28_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork15_outs_0,
      outs(1) => fork15_outs_1,
      outs(2) => fork15_outs_2,
      outs(3) => fork15_outs_3,
      outs(4) => fork15_outs_4,
      outs_valid(0) => fork15_outs_0_valid,
      outs_valid(1) => fork15_outs_1_valid,
      outs_valid(2) => fork15_outs_2_valid,
      outs_valid(3) => fork15_outs_3_valid,
      outs_valid(4) => fork15_outs_4_valid,
      outs_ready(0) => fork15_outs_0_ready,
      outs_ready(1) => fork15_outs_1_ready,
      outs_ready(2) => fork15_outs_2_ready,
      outs_ready(3) => fork15_outs_3_ready,
      outs_ready(4) => fork15_outs_4_ready
    );

  mux2 : entity work.mux(arch) generic map(2, 3, 1)
    port map(
      index => fork16_outs_0,
      index_valid => fork16_outs_0_valid,
      index_ready => fork16_outs_0_ready,
      ins(0) => buffer13_outs,
      ins(1) => cond_br4_trueOut,
      ins_valid(0) => buffer13_outs_valid,
      ins_valid(1) => cond_br4_trueOut_valid,
      ins_ready(0) => buffer13_outs_ready,
      ins_ready(1) => cond_br4_trueOut_ready,
      clk => clk,
      rst => rst,
      outs => mux2_outs,
      outs_valid => mux2_outs_valid,
      outs_ready => mux2_outs_ready
    );

  control_merge1 : entity work.control_merge_dataless(arch) generic map(2, 1)
    port map(
      ins_valid(0) => fork3_outs_1_valid,
      ins_valid(1) => cond_br5_trueOut_valid,
      ins_ready(0) => fork3_outs_1_ready,
      ins_ready(1) => cond_br5_trueOut_ready,
      clk => clk,
      rst => rst,
      outs_valid => control_merge1_outs_valid,
      outs_ready => control_merge1_outs_ready,
      index => control_merge1_index,
      index_valid => control_merge1_index_valid,
      index_ready => control_merge1_index_ready
    );

  fork16 : entity work.handshake_fork(arch) generic map(2, 1)
    port map(
      ins => control_merge1_index,
      ins_valid => control_merge1_index_valid,
      ins_ready => control_merge1_index_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork16_outs_0,
      outs(1) => fork16_outs_1,
      outs_valid(0) => fork16_outs_0_valid,
      outs_valid(1) => fork16_outs_1_valid,
      outs_ready(0) => fork16_outs_0_ready,
      outs_ready(1) => fork16_outs_1_ready
    );

  buffer36 : entity work.oehb_dataless(arch)
    port map(
      ins_valid => control_merge1_outs_valid,
      ins_ready => control_merge1_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer36_outs_valid,
      outs_ready => buffer36_outs_ready
    );

  fork17 : entity work.fork_dataless(arch) generic map(2)
    port map(
      ins_valid => buffer36_outs_valid,
      ins_ready => buffer36_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid(0) => fork17_outs_0_valid,
      outs_valid(1) => fork17_outs_1_valid,
      outs_ready(0) => fork17_outs_0_ready,
      outs_ready(1) => fork17_outs_1_ready
    );

  constant16 : entity work.handshake_constant_2(arch) generic map(2)
    port map(
      ctrl_valid => fork17_outs_0_valid,
      ctrl_ready => fork17_outs_0_ready,
      clk => clk,
      rst => rst,
      outs => constant16_outs,
      outs_valid => constant16_outs_valid,
      outs_ready => constant16_outs_ready
    );

  fork18 : entity work.handshake_fork(arch) generic map(4, 2)
    port map(
      ins => constant16_outs,
      ins_valid => constant16_outs_valid,
      ins_ready => constant16_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork18_outs_0,
      outs(1) => fork18_outs_1,
      outs(2) => fork18_outs_2,
      outs(3) => fork18_outs_3,
      outs_valid(0) => fork18_outs_0_valid,
      outs_valid(1) => fork18_outs_1_valid,
      outs_valid(2) => fork18_outs_2_valid,
      outs_valid(3) => fork18_outs_3_valid,
      outs_ready(0) => fork18_outs_0_ready,
      outs_ready(1) => fork18_outs_1_ready,
      outs_ready(2) => fork18_outs_2_ready,
      outs_ready(3) => fork18_outs_3_ready
    );

  extsi29 : entity work.extsi(arch) generic map(2, 9)
    port map(
      ins => fork18_outs_0,
      ins_valid => fork18_outs_0_valid,
      ins_ready => fork18_outs_0_ready,
      clk => clk,
      rst => rst,
      outs => extsi29_outs,
      outs_valid => extsi29_outs_valid,
      outs_ready => extsi29_outs_ready
    );

  extsi30 : entity work.extsi(arch) generic map(2, 9)
    port map(
      ins => fork18_outs_1,
      ins_valid => fork18_outs_1_valid,
      ins_ready => fork18_outs_1_ready,
      clk => clk,
      rst => rst,
      outs => extsi30_outs,
      outs_valid => extsi30_outs_valid,
      outs_ready => extsi30_outs_ready
    );

  extsi11 : entity work.extsi(arch) generic map(2, 32)
    port map(
      ins => fork18_outs_3,
      ins_valid => fork18_outs_3_valid,
      ins_ready => fork18_outs_3_ready,
      clk => clk,
      rst => rst,
      outs => extsi11_outs,
      outs_valid => extsi11_outs_valid,
      outs_ready => extsi11_outs_ready
    );

  source0 : entity work.source(arch)
    port map(
      clk => clk,
      rst => rst,
      outs_valid => source0_outs_valid,
      outs_ready => source0_outs_ready
    );

  constant7 : entity work.handshake_constant_3(arch) generic map(32)
    port map(
      ctrl_valid => source0_outs_valid,
      ctrl_ready => source0_outs_ready,
      clk => clk,
      rst => rst,
      outs => constant7_outs,
      outs_valid => constant7_outs_valid,
      outs_ready => constant7_outs_ready
    );

  source1 : entity work.source(arch)
    port map(
      clk => clk,
      rst => rst,
      outs_valid => source1_outs_valid,
      outs_ready => source1_outs_ready
    );

  constant18 : entity work.handshake_constant_4(arch) generic map(8)
    port map(
      ctrl_valid => source1_outs_valid,
      ctrl_ready => source1_outs_ready,
      clk => clk,
      rst => rst,
      outs => constant18_outs,
      outs_valid => constant18_outs_valid,
      outs_ready => constant18_outs_ready
    );

  extsi31 : entity work.extsi(arch) generic map(8, 9)
    port map(
      ins => constant18_outs,
      ins_valid => constant18_outs_valid,
      ins_ready => constant18_outs_ready,
      clk => clk,
      rst => rst,
      outs => extsi31_outs,
      outs_valid => extsi31_outs_valid,
      outs_ready => extsi31_outs_ready
    );

  source2 : entity work.source(arch)
    port map(
      clk => clk,
      rst => rst,
      outs_valid => source2_outs_valid,
      outs_ready => source2_outs_ready
    );

  constant19 : entity work.handshake_constant_2(arch) generic map(2)
    port map(
      ctrl_valid => source2_outs_valid,
      ctrl_ready => source2_outs_ready,
      clk => clk,
      rst => rst,
      outs => constant19_outs,
      outs_valid => constant19_outs_valid,
      outs_ready => constant19_outs_ready
    );

  extsi13 : entity work.extsi(arch) generic map(2, 32)
    port map(
      ins => constant19_outs,
      ins_valid => constant19_outs_valid,
      ins_ready => constant19_outs_ready,
      clk => clk,
      rst => rst,
      outs => extsi13_outs,
      outs_valid => extsi13_outs_valid,
      outs_ready => extsi13_outs_ready
    );

  addi2 : entity work.addi(arch) generic map(32)
    port map(
      lhs => fork15_outs_0,
      lhs_valid => fork15_outs_0_valid,
      lhs_ready => fork15_outs_0_ready,
      rhs => constant7_outs,
      rhs_valid => constant7_outs_valid,
      rhs_ready => constant7_outs_ready,
      clk => clk,
      rst => rst,
      result => addi2_result,
      result_valid => addi2_result_valid,
      result_ready => addi2_result_ready
    );

  buffer39 : entity work.oehb(arch) generic map(32)
    port map(
      ins => addi2_result,
      ins_valid => addi2_result_valid,
      ins_ready => addi2_result_ready,
      clk => clk,
      rst => rst,
      outs => buffer39_outs,
      outs_valid => buffer39_outs_valid,
      outs_ready => buffer39_outs_ready
    );

  fork19 : entity work.handshake_fork(arch) generic map(3, 32)
    port map(
      ins => buffer39_outs,
      ins_valid => buffer39_outs_valid,
      ins_ready => buffer39_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork19_outs_0,
      outs(1) => fork19_outs_1,
      outs(2) => fork19_outs_2,
      outs_valid(0) => fork19_outs_0_valid,
      outs_valid(1) => fork19_outs_1_valid,
      outs_valid(2) => fork19_outs_2_valid,
      outs_ready(0) => fork19_outs_0_ready,
      outs_ready(1) => fork19_outs_1_ready,
      outs_ready(2) => fork19_outs_2_ready
    );

  buffer0 : entity work.tfifo(arch) generic map(1, 32)
    port map(
      ins => fork19_outs_2,
      ins_valid => fork19_outs_2_valid,
      ins_ready => fork19_outs_2_ready,
      clk => clk,
      rst => rst,
      outs => buffer0_outs,
      outs_valid => buffer0_outs_valid,
      outs_ready => buffer0_outs_ready
    );

  fork20 : entity work.handshake_fork(arch) generic map(2, 32)
    port map(
      ins => buffer0_outs,
      ins_valid => buffer0_outs_valid,
      ins_ready => buffer0_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork20_outs_0,
      outs(1) => fork20_outs_1,
      outs_valid(0) => fork20_outs_0_valid,
      outs_valid(1) => fork20_outs_1_valid,
      outs_ready(0) => fork20_outs_0_ready,
      outs_ready(1) => fork20_outs_1_ready
    );

  init80 : entity work.tehb_init(arch) generic map(32, 0)
    port map(
      ins => fork20_outs_0,
      ins_valid => fork20_outs_0_valid,
      ins_ready => fork20_outs_0_ready,
      clk => clk,
      rst => rst,
      outs => init80_outs,
      outs_valid => init80_outs_valid,
      outs_ready => init80_outs_ready
    );

  buffer1 : entity work.tfifo_dataless(arch) generic map(1)
    port map(
      ins_valid => unbundle4_outs_0_valid,
      ins_ready => unbundle4_outs_0_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer1_outs_valid,
      outs_ready => buffer1_outs_ready
    );

  fork21 : entity work.fork_dataless(arch) generic map(2)
    port map(
      ins_valid => buffer1_outs_valid,
      ins_ready => buffer1_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid(0) => fork21_outs_0_valid,
      outs_valid(1) => fork21_outs_1_valid,
      outs_ready(0) => fork21_outs_0_ready,
      outs_ready(1) => fork21_outs_1_ready
    );

  init81 : entity work.tehb_dataless_init(arch)
    port map(
      ins_valid => fork21_outs_0_valid,
      ins_ready => fork21_outs_0_ready,
      clk => clk,
      rst => rst,
      outs_valid => init81_outs_valid,
      outs_ready => init81_outs_ready
    );

  fork22 : entity work.fork_dataless(arch) generic map(2)
    port map(
      ins_valid => init81_outs_valid,
      ins_ready => init81_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid(0) => fork22_outs_0_valid,
      outs_valid(1) => fork22_outs_1_valid,
      outs_ready(0) => fork22_outs_0_ready,
      outs_ready(1) => fork22_outs_1_ready
    );

  init82 : entity work.tehb_dataless_init(arch)
    port map(
      ins_valid => fork22_outs_0_valid,
      ins_ready => fork22_outs_0_ready,
      clk => clk,
      rst => rst,
      outs_valid => init82_outs_valid,
      outs_ready => init82_outs_ready
    );

  gate0 : entity work.gate(arch) generic map(2, 32)
    port map(
      ins(0) => fork19_outs_1,
      ins_valid(0) => fork19_outs_1_valid,
      ins_valid(1) => fork5_outs_11_valid,
      ins_ready(0) => fork19_outs_1_ready,
      ins_ready(1) => fork5_outs_11_ready,
      clk => clk,
      rst => rst,
      outs => gate0_outs,
      outs_valid => gate0_outs_valid,
      outs_ready => gate0_outs_ready
    );

  fork23 : entity work.handshake_fork(arch) generic map(2, 32)
    port map(
      ins => gate0_outs,
      ins_valid => gate0_outs_valid,
      ins_ready => gate0_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork23_outs_0,
      outs(1) => fork23_outs_1,
      outs_valid(0) => fork23_outs_0_valid,
      outs_valid(1) => fork23_outs_1_valid,
      outs_ready(0) => fork23_outs_0_ready,
      outs_ready(1) => fork23_outs_1_ready
    );

  cmpi3 : entity work.handshake_cmpi_0(arch) generic map(32)
    port map(
      lhs => fork23_outs_1,
      lhs_valid => fork23_outs_1_valid,
      lhs_ready => fork23_outs_1_ready,
      rhs => extsi23_outs,
      rhs_valid => extsi23_outs_valid,
      rhs_ready => extsi23_outs_ready,
      clk => clk,
      rst => rst,
      result => cmpi3_result,
      result_valid => cmpi3_result_valid,
      result_ready => cmpi3_result_ready
    );

  fork24 : entity work.handshake_fork(arch) generic map(2, 1)
    port map(
      ins => cmpi3_result,
      ins_valid => cmpi3_result_valid,
      ins_ready => cmpi3_result_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork24_outs_0,
      outs(1) => fork24_outs_1,
      outs_valid(0) => fork24_outs_0_valid,
      outs_valid(1) => fork24_outs_1_valid,
      outs_ready(0) => fork24_outs_0_ready,
      outs_ready(1) => fork24_outs_1_ready
    );

  cmpi4 : entity work.handshake_cmpi_0(arch) generic map(32)
    port map(
      lhs => fork23_outs_0,
      lhs_valid => fork23_outs_0_valid,
      lhs_ready => fork23_outs_0_ready,
      rhs => fork9_outs_0,
      rhs_valid => fork9_outs_0_valid,
      rhs_ready => fork9_outs_0_ready,
      clk => clk,
      rst => rst,
      result => cmpi4_result,
      result_valid => cmpi4_result_valid,
      result_ready => cmpi4_result_ready
    );

  fork25 : entity work.handshake_fork(arch) generic map(2, 1)
    port map(
      ins => cmpi4_result,
      ins_valid => cmpi4_result_valid,
      ins_ready => cmpi4_result_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork25_outs_0,
      outs(1) => fork25_outs_1,
      outs_valid(0) => fork25_outs_0_valid,
      outs_valid(1) => fork25_outs_1_valid,
      outs_ready(0) => fork25_outs_0_ready,
      outs_ready(1) => fork25_outs_1_ready
    );

  cond_br89 : entity work.cond_br_dataless(arch)
    port map(
      condition => fork24_outs_1,
      condition_valid => fork24_outs_1_valid,
      condition_ready => fork24_outs_1_ready,
      data_valid => fork5_outs_10_valid,
      data_ready => fork5_outs_10_ready,
      clk => clk,
      rst => rst,
      trueOut_valid => cond_br89_trueOut_valid,
      trueOut_ready => cond_br89_trueOut_ready,
      falseOut_valid => cond_br89_falseOut_valid,
      falseOut_ready => cond_br89_falseOut_ready
    );

  sink29 : entity work.sink_dataless(arch)
    port map(
      ins_valid => cond_br89_trueOut_valid,
      ins_ready => cond_br89_trueOut_ready,
      clk => clk,
      rst => rst
    );

  cond_br90 : entity work.cond_br_dataless(arch)
    port map(
      condition => fork25_outs_1,
      condition_valid => fork25_outs_1_valid,
      condition_ready => fork25_outs_1_ready,
      data_valid => fork5_outs_9_valid,
      data_ready => fork5_outs_9_ready,
      clk => clk,
      rst => rst,
      trueOut_valid => cond_br90_trueOut_valid,
      trueOut_ready => cond_br90_trueOut_ready,
      falseOut_valid => cond_br90_falseOut_valid,
      falseOut_ready => cond_br90_falseOut_ready
    );

  sink30 : entity work.sink_dataless(arch)
    port map(
      ins_valid => cond_br90_trueOut_valid,
      ins_ready => cond_br90_trueOut_ready,
      clk => clk,
      rst => rst
    );

  source7 : entity work.source(arch)
    port map(
      clk => clk,
      rst => rst,
      outs_valid => source7_outs_valid,
      outs_ready => source7_outs_ready
    );

  mux85 : entity work.mux_dataless(arch) generic map(2, 1)
    port map(
      index => fork24_outs_0,
      index_valid => fork24_outs_0_valid,
      index_ready => fork24_outs_0_ready,
      ins_valid(0) => cond_br89_falseOut_valid,
      ins_valid(1) => source7_outs_valid,
      ins_ready(0) => cond_br89_falseOut_ready,
      ins_ready(1) => source7_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => mux85_outs_valid,
      outs_ready => mux85_outs_ready
    );

  source8 : entity work.source(arch)
    port map(
      clk => clk,
      rst => rst,
      outs_valid => source8_outs_valid,
      outs_ready => source8_outs_ready
    );

  mux86 : entity work.mux_dataless(arch) generic map(2, 1)
    port map(
      index => fork25_outs_0,
      index_valid => fork25_outs_0_valid,
      index_ready => fork25_outs_0_ready,
      ins_valid(0) => cond_br90_falseOut_valid,
      ins_valid(1) => source8_outs_valid,
      ins_ready(0) => cond_br90_falseOut_ready,
      ins_ready(1) => source8_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => mux86_outs_valid,
      outs_ready => mux86_outs_ready
    );

  buffer40 : entity work.tehb_dataless(arch)
    port map(
      ins_valid => mux85_outs_valid,
      ins_ready => mux85_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer40_outs_valid,
      outs_ready => buffer40_outs_ready
    );

  buffer41 : entity work.tehb_dataless(arch)
    port map(
      ins_valid => mux86_outs_valid,
      ins_ready => mux86_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer41_outs_valid,
      outs_ready => buffer41_outs_ready
    );

  join0 : entity work.join_handshake(arch) generic map(2)
    port map(
      ins_valid(0) => buffer40_outs_valid,
      ins_valid(1) => buffer41_outs_valid,
      ins_ready(0) => buffer40_outs_ready,
      ins_ready(1) => buffer41_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => join0_outs_valid,
      outs_ready => join0_outs_ready
    );

  gate1 : entity work.gate(arch) generic map(2, 32)
    port map(
      ins(0) => fork19_outs_0,
      ins_valid(0) => fork19_outs_0_valid,
      ins_valid(1) => join0_outs_valid,
      ins_ready(0) => fork19_outs_0_ready,
      ins_ready(1) => join0_outs_ready,
      clk => clk,
      rst => rst,
      outs => gate1_outs,
      outs_valid => gate1_outs_valid,
      outs_ready => gate1_outs_ready
    );

  trunci0 : entity work.trunci(arch) generic map(32, 7)
    port map(
      ins => gate1_outs,
      ins_valid => gate1_outs_valid,
      ins_ready => gate1_outs_ready,
      clk => clk,
      rst => rst,
      outs => trunci0_outs,
      outs_valid => trunci0_outs_valid,
      outs_ready => trunci0_outs_ready
    );

  load0 : entity work.load(arch) generic map(32, 7)
    port map(
      addrIn => trunci0_outs,
      addrIn_valid => trunci0_outs_valid,
      addrIn_ready => trunci0_outs_ready,
      dataFromMem => mem_controller1_ldData_0,
      dataFromMem_valid => mem_controller1_ldData_0_valid,
      dataFromMem_ready => mem_controller1_ldData_0_ready,
      clk => clk,
      rst => rst,
      addrOut => load0_addrOut,
      addrOut_valid => load0_addrOut_valid,
      addrOut_ready => load0_addrOut_ready,
      dataOut => load0_dataOut,
      dataOut_valid => load0_dataOut_valid,
      dataOut_ready => load0_dataOut_ready
    );

  fork26 : entity work.handshake_fork(arch) generic map(2, 32)
    port map(
      ins => load0_dataOut,
      ins_valid => load0_dataOut_valid,
      ins_ready => load0_dataOut_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork26_outs_0,
      outs(1) => fork26_outs_1,
      outs_valid(0) => fork26_outs_0_valid,
      outs_valid(1) => fork26_outs_1_valid,
      outs_ready(0) => fork26_outs_0_ready,
      outs_ready(1) => fork26_outs_1_ready
    );

  buffer2 : entity work.tfifo(arch) generic map(1, 8)
    port map(
      ins => fork14_outs_3,
      ins_valid => fork14_outs_3_valid,
      ins_ready => fork14_outs_3_ready,
      clk => clk,
      rst => rst,
      outs => buffer2_outs,
      outs_valid => buffer2_outs_valid,
      outs_ready => buffer2_outs_ready
    );

  fork27 : entity work.handshake_fork(arch) generic map(2, 8)
    port map(
      ins => buffer2_outs,
      ins_valid => buffer2_outs_valid,
      ins_ready => buffer2_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork27_outs_0,
      outs(1) => fork27_outs_1,
      outs_valid(0) => fork27_outs_0_valid,
      outs_valid(1) => fork27_outs_1_valid,
      outs_ready(0) => fork27_outs_0_ready,
      outs_ready(1) => fork27_outs_1_ready
    );

  extsi32 : entity work.extsi(arch) generic map(8, 32)
    port map(
      ins => fork27_outs_1,
      ins_valid => fork27_outs_1_valid,
      ins_ready => fork27_outs_1_ready,
      clk => clk,
      rst => rst,
      outs => extsi32_outs,
      outs_valid => extsi32_outs_valid,
      outs_ready => extsi32_outs_ready
    );

  init83 : entity work.tehb_init(arch) generic map(32, 0)
    port map(
      ins => extsi32_outs,
      ins_valid => extsi32_outs_valid,
      ins_ready => extsi32_outs_ready,
      clk => clk,
      rst => rst,
      outs => init83_outs,
      outs_valid => init83_outs_valid,
      outs_ready => init83_outs_ready
    );

  buffer3 : entity work.tfifo_dataless(arch) generic map(1)
    port map(
      ins_valid => unbundle3_outs_0_valid,
      ins_ready => unbundle3_outs_0_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer3_outs_valid,
      outs_ready => buffer3_outs_ready
    );

  fork28 : entity work.fork_dataless(arch) generic map(2)
    port map(
      ins_valid => buffer3_outs_valid,
      ins_ready => buffer3_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid(0) => fork28_outs_0_valid,
      outs_valid(1) => fork28_outs_1_valid,
      outs_ready(0) => fork28_outs_0_ready,
      outs_ready(1) => fork28_outs_1_ready
    );

  init84 : entity work.tehb_dataless_init(arch)
    port map(
      ins_valid => fork28_outs_0_valid,
      ins_ready => fork28_outs_0_ready,
      clk => clk,
      rst => rst,
      outs_valid => init84_outs_valid,
      outs_ready => init84_outs_ready
    );

  fork29 : entity work.fork_dataless(arch) generic map(2)
    port map(
      ins_valid => init84_outs_valid,
      ins_ready => init84_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid(0) => fork29_outs_0_valid,
      outs_valid(1) => fork29_outs_1_valid,
      outs_ready(0) => fork29_outs_0_ready,
      outs_ready(1) => fork29_outs_1_ready
    );

  init85 : entity work.tehb_dataless_init(arch)
    port map(
      ins_valid => fork29_outs_0_valid,
      ins_ready => fork29_outs_0_ready,
      clk => clk,
      rst => rst,
      outs_valid => init85_outs_valid,
      outs_ready => init85_outs_ready
    );

  gate2 : entity work.gate(arch) generic map(2, 32)
    port map(
      ins(0) => fork15_outs_1,
      ins_valid(0) => fork15_outs_1_valid,
      ins_valid(1) => fork5_outs_8_valid,
      ins_ready(0) => fork15_outs_1_ready,
      ins_ready(1) => fork5_outs_8_ready,
      clk => clk,
      rst => rst,
      outs => gate2_outs,
      outs_valid => gate2_outs_valid,
      outs_ready => gate2_outs_ready
    );

  fork30 : entity work.handshake_fork(arch) generic map(2, 32)
    port map(
      ins => gate2_outs,
      ins_valid => gate2_outs_valid,
      ins_ready => gate2_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork30_outs_0,
      outs(1) => fork30_outs_1,
      outs_valid(0) => fork30_outs_0_valid,
      outs_valid(1) => fork30_outs_1_valid,
      outs_ready(0) => fork30_outs_0_ready,
      outs_ready(1) => fork30_outs_1_ready
    );

  cmpi5 : entity work.handshake_cmpi_0(arch) generic map(32)
    port map(
      lhs => fork30_outs_1,
      lhs_valid => fork30_outs_1_valid,
      lhs_ready => fork30_outs_1_ready,
      rhs => extsi22_outs,
      rhs_valid => extsi22_outs_valid,
      rhs_ready => extsi22_outs_ready,
      clk => clk,
      rst => rst,
      result => cmpi5_result,
      result_valid => cmpi5_result_valid,
      result_ready => cmpi5_result_ready
    );

  fork31 : entity work.handshake_fork(arch) generic map(2, 1)
    port map(
      ins => cmpi5_result,
      ins_valid => cmpi5_result_valid,
      ins_ready => cmpi5_result_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork31_outs_0,
      outs(1) => fork31_outs_1,
      outs_valid(0) => fork31_outs_0_valid,
      outs_valid(1) => fork31_outs_1_valid,
      outs_ready(0) => fork31_outs_0_ready,
      outs_ready(1) => fork31_outs_1_ready
    );

  cmpi6 : entity work.handshake_cmpi_0(arch) generic map(32)
    port map(
      lhs => fork30_outs_0,
      lhs_valid => fork30_outs_0_valid,
      lhs_ready => fork30_outs_0_ready,
      rhs => fork6_outs_0,
      rhs_valid => fork6_outs_0_valid,
      rhs_ready => fork6_outs_0_ready,
      clk => clk,
      rst => rst,
      result => cmpi6_result,
      result_valid => cmpi6_result_valid,
      result_ready => cmpi6_result_ready
    );

  fork32 : entity work.handshake_fork(arch) generic map(2, 1)
    port map(
      ins => cmpi6_result,
      ins_valid => cmpi6_result_valid,
      ins_ready => cmpi6_result_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork32_outs_0,
      outs(1) => fork32_outs_1,
      outs_valid(0) => fork32_outs_0_valid,
      outs_valid(1) => fork32_outs_1_valid,
      outs_ready(0) => fork32_outs_0_ready,
      outs_ready(1) => fork32_outs_1_ready
    );

  cond_br91 : entity work.cond_br_dataless(arch)
    port map(
      condition => fork31_outs_1,
      condition_valid => fork31_outs_1_valid,
      condition_ready => fork31_outs_1_ready,
      data_valid => fork5_outs_7_valid,
      data_ready => fork5_outs_7_ready,
      clk => clk,
      rst => rst,
      trueOut_valid => cond_br91_trueOut_valid,
      trueOut_ready => cond_br91_trueOut_ready,
      falseOut_valid => cond_br91_falseOut_valid,
      falseOut_ready => cond_br91_falseOut_ready
    );

  sink31 : entity work.sink_dataless(arch)
    port map(
      ins_valid => cond_br91_trueOut_valid,
      ins_ready => cond_br91_trueOut_ready,
      clk => clk,
      rst => rst
    );

  cond_br92 : entity work.cond_br_dataless(arch)
    port map(
      condition => fork32_outs_1,
      condition_valid => fork32_outs_1_valid,
      condition_ready => fork32_outs_1_ready,
      data_valid => fork5_outs_6_valid,
      data_ready => fork5_outs_6_ready,
      clk => clk,
      rst => rst,
      trueOut_valid => cond_br92_trueOut_valid,
      trueOut_ready => cond_br92_trueOut_ready,
      falseOut_valid => cond_br92_falseOut_valid,
      falseOut_ready => cond_br92_falseOut_ready
    );

  sink32 : entity work.sink_dataless(arch)
    port map(
      ins_valid => cond_br92_trueOut_valid,
      ins_ready => cond_br92_trueOut_ready,
      clk => clk,
      rst => rst
    );

  source9 : entity work.source(arch)
    port map(
      clk => clk,
      rst => rst,
      outs_valid => source9_outs_valid,
      outs_ready => source9_outs_ready
    );

  mux87 : entity work.mux_dataless(arch) generic map(2, 1)
    port map(
      index => fork31_outs_0,
      index_valid => fork31_outs_0_valid,
      index_ready => fork31_outs_0_ready,
      ins_valid(0) => cond_br91_falseOut_valid,
      ins_valid(1) => source9_outs_valid,
      ins_ready(0) => cond_br91_falseOut_ready,
      ins_ready(1) => source9_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => mux87_outs_valid,
      outs_ready => mux87_outs_ready
    );

  source10 : entity work.source(arch)
    port map(
      clk => clk,
      rst => rst,
      outs_valid => source10_outs_valid,
      outs_ready => source10_outs_ready
    );

  mux88 : entity work.mux_dataless(arch) generic map(2, 1)
    port map(
      index => fork32_outs_0,
      index_valid => fork32_outs_0_valid,
      index_ready => fork32_outs_0_ready,
      ins_valid(0) => cond_br92_falseOut_valid,
      ins_valid(1) => source10_outs_valid,
      ins_ready(0) => cond_br92_falseOut_ready,
      ins_ready(1) => source10_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => mux88_outs_valid,
      outs_ready => mux88_outs_ready
    );

  buffer42 : entity work.tehb_dataless(arch)
    port map(
      ins_valid => mux87_outs_valid,
      ins_ready => mux87_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer42_outs_valid,
      outs_ready => buffer42_outs_ready
    );

  buffer43 : entity work.tehb_dataless(arch)
    port map(
      ins_valid => mux88_outs_valid,
      ins_ready => mux88_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer43_outs_valid,
      outs_ready => buffer43_outs_ready
    );

  join1 : entity work.join_handshake(arch) generic map(2)
    port map(
      ins_valid(0) => buffer42_outs_valid,
      ins_valid(1) => buffer43_outs_valid,
      ins_ready(0) => buffer42_outs_ready,
      ins_ready(1) => buffer43_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => join1_outs_valid,
      outs_ready => join1_outs_ready
    );

  gate3 : entity work.gate(arch) generic map(2, 32)
    port map(
      ins(0) => fork15_outs_2,
      ins_valid(0) => fork15_outs_2_valid,
      ins_valid(1) => join1_outs_valid,
      ins_ready(0) => fork15_outs_2_ready,
      ins_ready(1) => join1_outs_ready,
      clk => clk,
      rst => rst,
      outs => gate3_outs,
      outs_valid => gate3_outs_valid,
      outs_ready => gate3_outs_ready
    );

  trunci1 : entity work.trunci(arch) generic map(32, 7)
    port map(
      ins => gate3_outs,
      ins_valid => gate3_outs_valid,
      ins_ready => gate3_outs_ready,
      clk => clk,
      rst => rst,
      outs => trunci1_outs,
      outs_valid => trunci1_outs_valid,
      outs_ready => trunci1_outs_ready
    );

  load1 : entity work.load(arch) generic map(32, 7)
    port map(
      addrIn => trunci1_outs,
      addrIn_valid => trunci1_outs_valid,
      addrIn_ready => trunci1_outs_ready,
      dataFromMem => mem_controller1_ldData_1,
      dataFromMem_valid => mem_controller1_ldData_1_valid,
      dataFromMem_ready => mem_controller1_ldData_1_ready,
      clk => clk,
      rst => rst,
      addrOut => load1_addrOut,
      addrOut_valid => load1_addrOut_valid,
      addrOut_ready => load1_addrOut_ready,
      dataOut => load1_dataOut,
      dataOut_valid => load1_dataOut_valid,
      dataOut_ready => load1_dataOut_ready
    );

  fork33 : entity work.handshake_fork(arch) generic map(2, 32)
    port map(
      ins => load1_dataOut,
      ins_valid => load1_dataOut_valid,
      ins_ready => load1_dataOut_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork33_outs_0,
      outs(1) => fork33_outs_1,
      outs_valid(0) => fork33_outs_0_valid,
      outs_valid(1) => fork33_outs_1_valid,
      outs_ready(0) => fork33_outs_0_ready,
      outs_ready(1) => fork33_outs_1_ready
    );

  addi0 : entity work.addi(arch) generic map(32)
    port map(
      lhs => fork26_outs_1,
      lhs_valid => fork26_outs_1_valid,
      lhs_ready => fork26_outs_1_ready,
      rhs => fork33_outs_1,
      rhs_valid => fork33_outs_1_valid,
      rhs_ready => fork33_outs_1_ready,
      clk => clk,
      rst => rst,
      result => addi0_result,
      result_valid => addi0_result_valid,
      result_ready => addi0_result_ready
    );

  addi3 : entity work.addi(arch) generic map(9)
    port map(
      lhs => extsi27_outs,
      lhs_valid => extsi27_outs_valid,
      lhs_ready => extsi27_outs_ready,
      rhs => extsi30_outs,
      rhs_valid => extsi30_outs_valid,
      rhs_ready => extsi30_outs_ready,
      clk => clk,
      rst => rst,
      result => addi3_result,
      result_valid => addi3_result_valid,
      result_ready => addi3_result_ready
    );

  buffer45 : entity work.oehb(arch) generic map(9)
    port map(
      ins => addi3_result,
      ins_valid => addi3_result_valid,
      ins_ready => addi3_result_ready,
      clk => clk,
      rst => rst,
      outs => buffer45_outs,
      outs_valid => buffer45_outs_valid,
      outs_ready => buffer45_outs_ready
    );

  fork34 : entity work.handshake_fork(arch) generic map(2, 9)
    port map(
      ins => buffer45_outs,
      ins_valid => buffer45_outs_valid,
      ins_ready => buffer45_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork34_outs_0,
      outs(1) => fork34_outs_1,
      outs_valid(0) => fork34_outs_0_valid,
      outs_valid(1) => fork34_outs_1_valid,
      outs_ready(0) => fork34_outs_0_ready,
      outs_ready(1) => fork34_outs_1_ready
    );

  extsi33 : entity work.extsi(arch) generic map(9, 32)
    port map(
      ins => buffer123_outs,
      ins_valid => buffer123_outs_valid,
      ins_ready => buffer123_outs_ready,
      clk => clk,
      rst => rst,
      outs => extsi33_outs,
      outs_valid => extsi33_outs_valid,
      outs_ready => extsi33_outs_ready
    );

  buffer123 : entity work.tfifo(arch) generic map(1, 9)
    port map(
      ins => fork34_outs_1,
      ins_valid => fork34_outs_1_valid,
      ins_ready => fork34_outs_1_ready,
      clk => clk,
      rst => rst,
      outs => buffer123_outs,
      outs_valid => buffer123_outs_valid,
      outs_ready => buffer123_outs_ready
    );

  fork35 : entity work.handshake_fork(arch) generic map(2, 32)
    port map(
      ins => extsi33_outs,
      ins_valid => extsi33_outs_valid,
      ins_ready => extsi33_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork35_outs_0,
      outs(1) => fork35_outs_1,
      outs_valid(0) => fork35_outs_0_valid,
      outs_valid(1) => fork35_outs_1_valid,
      outs_ready(0) => fork35_outs_0_ready,
      outs_ready(1) => fork35_outs_1_ready
    );

  buffer4 : entity work.tfifo(arch) generic map(1, 9)
    port map(
      ins => fork34_outs_0,
      ins_valid => fork34_outs_0_valid,
      ins_ready => fork34_outs_0_ready,
      clk => clk,
      rst => rst,
      outs => buffer4_outs,
      outs_valid => buffer4_outs_valid,
      outs_ready => buffer4_outs_ready
    );

  fork36 : entity work.handshake_fork(arch) generic map(2, 9)
    port map(
      ins => buffer4_outs,
      ins_valid => buffer4_outs_valid,
      ins_ready => buffer4_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork36_outs_0,
      outs(1) => fork36_outs_1,
      outs_valid(0) => fork36_outs_0_valid,
      outs_valid(1) => fork36_outs_1_valid,
      outs_ready(0) => fork36_outs_0_ready,
      outs_ready(1) => fork36_outs_1_ready
    );

  extsi34 : entity work.extsi(arch) generic map(9, 32)
    port map(
      ins => fork36_outs_1,
      ins_valid => fork36_outs_1_valid,
      ins_ready => fork36_outs_1_ready,
      clk => clk,
      rst => rst,
      outs => extsi34_outs,
      outs_valid => extsi34_outs_valid,
      outs_ready => extsi34_outs_ready
    );

  init86 : entity work.tehb_init(arch) generic map(32, 0)
    port map(
      ins => extsi34_outs,
      ins_valid => extsi34_outs_valid,
      ins_ready => extsi34_outs_ready,
      clk => clk,
      rst => rst,
      outs => init86_outs,
      outs_valid => init86_outs_valid,
      outs_ready => init86_outs_ready
    );

  buffer5 : entity work.tfifo_dataless(arch) generic map(1)
    port map(
      ins_valid => unbundle5_outs_0_valid,
      ins_ready => unbundle5_outs_0_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer5_outs_valid,
      outs_ready => buffer5_outs_ready
    );

  fork37 : entity work.fork_dataless(arch) generic map(2)
    port map(
      ins_valid => buffer5_outs_valid,
      ins_ready => buffer5_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid(0) => fork37_outs_0_valid,
      outs_valid(1) => fork37_outs_1_valid,
      outs_ready(0) => fork37_outs_0_ready,
      outs_ready(1) => fork37_outs_1_ready
    );

  init87 : entity work.tehb_dataless_init(arch)
    port map(
      ins_valid => fork37_outs_0_valid,
      ins_ready => fork37_outs_0_ready,
      clk => clk,
      rst => rst,
      outs_valid => init87_outs_valid,
      outs_ready => init87_outs_ready
    );

  fork38 : entity work.fork_dataless(arch) generic map(2)
    port map(
      ins_valid => init87_outs_valid,
      ins_ready => init87_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid(0) => fork38_outs_0_valid,
      outs_valid(1) => fork38_outs_1_valid,
      outs_ready(0) => fork38_outs_0_ready,
      outs_ready(1) => fork38_outs_1_ready
    );

  init88 : entity work.tehb_dataless_init(arch)
    port map(
      ins_valid => fork38_outs_0_valid,
      ins_ready => fork38_outs_0_ready,
      clk => clk,
      rst => rst,
      outs_valid => init88_outs_valid,
      outs_ready => init88_outs_ready
    );

  gate4 : entity work.gate(arch) generic map(2, 32)
    port map(
      ins(0) => fork35_outs_0,
      ins_valid(0) => fork35_outs_0_valid,
      ins_valid(1) => fork5_outs_5_valid,
      ins_ready(0) => fork35_outs_0_ready,
      ins_ready(1) => fork5_outs_5_ready,
      clk => clk,
      rst => rst,
      outs => gate4_outs,
      outs_valid => gate4_outs_valid,
      outs_ready => gate4_outs_ready
    );

  fork39 : entity work.handshake_fork(arch) generic map(2, 32)
    port map(
      ins => gate4_outs,
      ins_valid => gate4_outs_valid,
      ins_ready => gate4_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork39_outs_0,
      outs(1) => fork39_outs_1,
      outs_valid(0) => fork39_outs_0_valid,
      outs_valid(1) => fork39_outs_1_valid,
      outs_ready(0) => fork39_outs_0_ready,
      outs_ready(1) => fork39_outs_1_ready
    );

  cmpi7 : entity work.handshake_cmpi_0(arch) generic map(32)
    port map(
      lhs => fork39_outs_1,
      lhs_valid => fork39_outs_1_valid,
      lhs_ready => fork39_outs_1_ready,
      rhs => extsi24_outs,
      rhs_valid => extsi24_outs_valid,
      rhs_ready => extsi24_outs_ready,
      clk => clk,
      rst => rst,
      result => cmpi7_result,
      result_valid => cmpi7_result_valid,
      result_ready => cmpi7_result_ready
    );

  fork40 : entity work.handshake_fork(arch) generic map(2, 1)
    port map(
      ins => cmpi7_result,
      ins_valid => cmpi7_result_valid,
      ins_ready => cmpi7_result_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork40_outs_0,
      outs(1) => fork40_outs_1,
      outs_valid(0) => fork40_outs_0_valid,
      outs_valid(1) => fork40_outs_1_valid,
      outs_ready(0) => fork40_outs_0_ready,
      outs_ready(1) => fork40_outs_1_ready
    );

  cmpi8 : entity work.handshake_cmpi_0(arch) generic map(32)
    port map(
      lhs => fork39_outs_0,
      lhs_valid => fork39_outs_0_valid,
      lhs_ready => fork39_outs_0_ready,
      rhs => fork10_outs_0,
      rhs_valid => fork10_outs_0_valid,
      rhs_ready => fork10_outs_0_ready,
      clk => clk,
      rst => rst,
      result => cmpi8_result,
      result_valid => cmpi8_result_valid,
      result_ready => cmpi8_result_ready
    );

  fork41 : entity work.handshake_fork(arch) generic map(2, 1)
    port map(
      ins => cmpi8_result,
      ins_valid => cmpi8_result_valid,
      ins_ready => cmpi8_result_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork41_outs_0,
      outs(1) => fork41_outs_1,
      outs_valid(0) => fork41_outs_0_valid,
      outs_valid(1) => fork41_outs_1_valid,
      outs_ready(0) => fork41_outs_0_ready,
      outs_ready(1) => fork41_outs_1_ready
    );

  cond_br93 : entity work.cond_br_dataless(arch)
    port map(
      condition => fork40_outs_1,
      condition_valid => fork40_outs_1_valid,
      condition_ready => fork40_outs_1_ready,
      data_valid => fork5_outs_4_valid,
      data_ready => fork5_outs_4_ready,
      clk => clk,
      rst => rst,
      trueOut_valid => cond_br93_trueOut_valid,
      trueOut_ready => cond_br93_trueOut_ready,
      falseOut_valid => cond_br93_falseOut_valid,
      falseOut_ready => cond_br93_falseOut_ready
    );

  sink33 : entity work.sink_dataless(arch)
    port map(
      ins_valid => cond_br93_trueOut_valid,
      ins_ready => cond_br93_trueOut_ready,
      clk => clk,
      rst => rst
    );

  cond_br94 : entity work.cond_br_dataless(arch)
    port map(
      condition => fork41_outs_1,
      condition_valid => fork41_outs_1_valid,
      condition_ready => fork41_outs_1_ready,
      data_valid => fork5_outs_3_valid,
      data_ready => fork5_outs_3_ready,
      clk => clk,
      rst => rst,
      trueOut_valid => cond_br94_trueOut_valid,
      trueOut_ready => cond_br94_trueOut_ready,
      falseOut_valid => cond_br94_falseOut_valid,
      falseOut_ready => cond_br94_falseOut_ready
    );

  sink34 : entity work.sink_dataless(arch)
    port map(
      ins_valid => cond_br94_trueOut_valid,
      ins_ready => cond_br94_trueOut_ready,
      clk => clk,
      rst => rst
    );

  source11 : entity work.source(arch)
    port map(
      clk => clk,
      rst => rst,
      outs_valid => source11_outs_valid,
      outs_ready => source11_outs_ready
    );

  mux89 : entity work.mux_dataless(arch) generic map(2, 1)
    port map(
      index => fork40_outs_0,
      index_valid => fork40_outs_0_valid,
      index_ready => fork40_outs_0_ready,
      ins_valid(0) => cond_br93_falseOut_valid,
      ins_valid(1) => source11_outs_valid,
      ins_ready(0) => cond_br93_falseOut_ready,
      ins_ready(1) => source11_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => mux89_outs_valid,
      outs_ready => mux89_outs_ready
    );

  source12 : entity work.source(arch)
    port map(
      clk => clk,
      rst => rst,
      outs_valid => source12_outs_valid,
      outs_ready => source12_outs_ready
    );

  mux90 : entity work.mux_dataless(arch) generic map(2, 1)
    port map(
      index => fork41_outs_0,
      index_valid => fork41_outs_0_valid,
      index_ready => fork41_outs_0_ready,
      ins_valid(0) => cond_br94_falseOut_valid,
      ins_valid(1) => source12_outs_valid,
      ins_ready(0) => cond_br94_falseOut_ready,
      ins_ready(1) => source12_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => mux90_outs_valid,
      outs_ready => mux90_outs_ready
    );

  buffer46 : entity work.tehb_dataless(arch)
    port map(
      ins_valid => mux89_outs_valid,
      ins_ready => mux89_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer46_outs_valid,
      outs_ready => buffer46_outs_ready
    );

  buffer47 : entity work.tehb_dataless(arch)
    port map(
      ins_valid => mux90_outs_valid,
      ins_ready => mux90_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer47_outs_valid,
      outs_ready => buffer47_outs_ready
    );

  join2 : entity work.join_handshake(arch) generic map(2)
    port map(
      ins_valid(0) => buffer46_outs_valid,
      ins_valid(1) => buffer47_outs_valid,
      ins_ready(0) => buffer46_outs_ready,
      ins_ready(1) => buffer47_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => join2_outs_valid,
      outs_ready => join2_outs_ready
    );

  gate5 : entity work.gate(arch) generic map(2, 32)
    port map(
      ins(0) => buffer134_outs,
      ins_valid(0) => buffer134_outs_valid,
      ins_valid(1) => join2_outs_valid,
      ins_ready(0) => buffer134_outs_ready,
      ins_ready(1) => join2_outs_ready,
      clk => clk,
      rst => rst,
      outs => gate5_outs,
      outs_valid => gate5_outs_valid,
      outs_ready => gate5_outs_ready
    );

  buffer134 : entity work.tfifo(arch) generic map(1, 32)
    port map(
      ins => fork35_outs_1,
      ins_valid => fork35_outs_1_valid,
      ins_ready => fork35_outs_1_ready,
      clk => clk,
      rst => rst,
      outs => buffer134_outs,
      outs_valid => buffer134_outs_valid,
      outs_ready => buffer134_outs_ready
    );

  trunci2 : entity work.trunci(arch) generic map(32, 7)
    port map(
      ins => gate5_outs,
      ins_valid => gate5_outs_valid,
      ins_ready => gate5_outs_ready,
      clk => clk,
      rst => rst,
      outs => trunci2_outs,
      outs_valid => trunci2_outs_valid,
      outs_ready => trunci2_outs_ready
    );

  load2 : entity work.load(arch) generic map(32, 7)
    port map(
      addrIn => trunci2_outs,
      addrIn_valid => trunci2_outs_valid,
      addrIn_ready => trunci2_outs_ready,
      dataFromMem => mem_controller1_ldData_2,
      dataFromMem_valid => mem_controller1_ldData_2_valid,
      dataFromMem_ready => mem_controller1_ldData_2_ready,
      clk => clk,
      rst => rst,
      addrOut => load2_addrOut,
      addrOut_valid => load2_addrOut_valid,
      addrOut_ready => load2_addrOut_ready,
      dataOut => load2_dataOut,
      dataOut_valid => load2_dataOut_valid,
      dataOut_ready => load2_dataOut_ready
    );

  fork42 : entity work.handshake_fork(arch) generic map(2, 32)
    port map(
      ins => load2_dataOut,
      ins_valid => load2_dataOut_valid,
      ins_ready => load2_dataOut_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork42_outs_0,
      outs(1) => fork42_outs_1,
      outs_valid(0) => fork42_outs_0_valid,
      outs_valid(1) => fork42_outs_1_valid,
      outs_ready(0) => fork42_outs_0_ready,
      outs_ready(1) => fork42_outs_1_ready
    );

  buffer44 : entity work.oehb(arch) generic map(32)
    port map(
      ins => addi0_result,
      ins_valid => addi0_result_valid,
      ins_ready => addi0_result_ready,
      clk => clk,
      rst => rst,
      outs => buffer44_outs,
      outs_valid => buffer44_outs_valid,
      outs_ready => buffer44_outs_ready
    );

  addi1 : entity work.addi(arch) generic map(32)
    port map(
      lhs => buffer44_outs,
      lhs_valid => buffer44_outs_valid,
      lhs_ready => buffer44_outs_ready,
      rhs => fork42_outs_1,
      rhs_valid => fork42_outs_1_valid,
      rhs_ready => fork42_outs_1_ready,
      clk => clk,
      rst => rst,
      result => addi1_result,
      result_valid => addi1_result_valid,
      result_ready => addi1_result_ready
    );

  buffer48 : entity work.oehb(arch) generic map(32)
    port map(
      ins => addi1_result,
      ins_valid => addi1_result_valid,
      ins_ready => addi1_result_ready,
      clk => clk,
      rst => rst,
      outs => buffer48_outs,
      outs_valid => buffer48_outs_valid,
      outs_ready => buffer48_outs_ready
    );

  fork43 : entity work.handshake_fork(arch) generic map(2, 32)
    port map(
      ins => buffer48_outs,
      ins_valid => buffer48_outs_valid,
      ins_ready => buffer48_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork43_outs_0,
      outs(1) => fork43_outs_1,
      outs_valid(0) => fork43_outs_0_valid,
      outs_valid(1) => fork43_outs_1_valid,
      outs_ready(0) => fork43_outs_0_ready,
      outs_ready(1) => fork43_outs_1_ready
    );

  shli0 : entity work.shli(arch) generic map(32)
    port map(
      lhs => fork43_outs_1,
      lhs_valid => fork43_outs_1_valid,
      lhs_ready => fork43_outs_1_ready,
      rhs => extsi13_outs,
      rhs_valid => extsi13_outs_valid,
      rhs_ready => extsi13_outs_ready,
      clk => clk,
      rst => rst,
      result => shli0_result,
      result_valid => shli0_result_valid,
      result_ready => shli0_result_ready
    );

  buffer49 : entity work.oehb(arch) generic map(32)
    port map(
      ins => shli0_result,
      ins_valid => shli0_result_valid,
      ins_ready => shli0_result_ready,
      clk => clk,
      rst => rst,
      outs => buffer49_outs,
      outs_valid => buffer49_outs_valid,
      outs_ready => buffer49_outs_ready
    );

  addi7 : entity work.addi(arch) generic map(32)
    port map(
      lhs => fork43_outs_0,
      lhs_valid => fork43_outs_0_valid,
      lhs_ready => fork43_outs_0_ready,
      rhs => buffer49_outs,
      rhs_valid => buffer49_outs_valid,
      rhs_ready => buffer49_outs_ready,
      clk => clk,
      rst => rst,
      result => addi7_result,
      result_valid => addi7_result_valid,
      result_ready => addi7_result_ready
    );

  buffer6 : entity work.tfifo(arch) generic map(1, 8)
    port map(
      ins => fork14_outs_1,
      ins_valid => fork14_outs_1_valid,
      ins_ready => fork14_outs_1_ready,
      clk => clk,
      rst => rst,
      outs => buffer6_outs,
      outs_valid => buffer6_outs_valid,
      outs_ready => buffer6_outs_ready
    );

  fork44 : entity work.handshake_fork(arch) generic map(2, 8)
    port map(
      ins => buffer6_outs,
      ins_valid => buffer6_outs_valid,
      ins_ready => buffer6_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork44_outs_0,
      outs(1) => fork44_outs_1,
      outs_valid(0) => fork44_outs_0_valid,
      outs_valid(1) => fork44_outs_1_valid,
      outs_ready(0) => fork44_outs_0_ready,
      outs_ready(1) => fork44_outs_1_ready
    );

  extsi35 : entity work.extsi(arch) generic map(8, 32)
    port map(
      ins => fork44_outs_1,
      ins_valid => fork44_outs_1_valid,
      ins_ready => fork44_outs_1_ready,
      clk => clk,
      rst => rst,
      outs => extsi35_outs,
      outs_valid => extsi35_outs_valid,
      outs_ready => extsi35_outs_ready
    );

  init89 : entity work.tehb_init(arch) generic map(32, 0)
    port map(
      ins => extsi35_outs,
      ins_valid => extsi35_outs_valid,
      ins_ready => extsi35_outs_ready,
      clk => clk,
      rst => rst,
      outs => init89_outs,
      outs_valid => init89_outs_valid,
      outs_ready => init89_outs_ready
    );

  buffer53 : entity work.oehb_dataless(arch)
    port map(
      ins_valid => store0_doneOut_valid,
      ins_ready => store0_doneOut_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer53_outs_valid,
      outs_ready => buffer53_outs_ready
    );

  buffer7 : entity work.tfifo_dataless(arch) generic map(1)
    port map(
      ins_valid => buffer53_outs_valid,
      ins_ready => buffer53_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer7_outs_valid,
      outs_ready => buffer7_outs_ready
    );

  fork45 : entity work.fork_dataless(arch) generic map(2)
    port map(
      ins_valid => buffer7_outs_valid,
      ins_ready => buffer7_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid(0) => fork45_outs_0_valid,
      outs_valid(1) => fork45_outs_1_valid,
      outs_ready(0) => fork45_outs_0_ready,
      outs_ready(1) => fork45_outs_1_ready
    );

  init90 : entity work.tehb_dataless_init(arch)
    port map(
      ins_valid => fork45_outs_0_valid,
      ins_ready => fork45_outs_0_ready,
      clk => clk,
      rst => rst,
      outs_valid => init90_outs_valid,
      outs_ready => init90_outs_ready
    );

  fork46 : entity work.fork_dataless(arch) generic map(2)
    port map(
      ins_valid => init90_outs_valid,
      ins_ready => init90_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid(0) => fork46_outs_0_valid,
      outs_valid(1) => fork46_outs_1_valid,
      outs_ready(0) => fork46_outs_0_ready,
      outs_ready(1) => fork46_outs_1_ready
    );

  init91 : entity work.tehb_dataless_init(arch)
    port map(
      ins_valid => fork46_outs_0_valid,
      ins_ready => fork46_outs_0_ready,
      clk => clk,
      rst => rst,
      outs_valid => init91_outs_valid,
      outs_ready => init91_outs_ready
    );

  gate6 : entity work.gate(arch) generic map(2, 32)
    port map(
      ins(0) => fork15_outs_3,
      ins_valid(0) => fork15_outs_3_valid,
      ins_valid(1) => fork5_outs_2_valid,
      ins_ready(0) => fork15_outs_3_ready,
      ins_ready(1) => fork5_outs_2_ready,
      clk => clk,
      rst => rst,
      outs => gate6_outs,
      outs_valid => gate6_outs_valid,
      outs_ready => gate6_outs_ready
    );

  fork47 : entity work.handshake_fork(arch) generic map(2, 32)
    port map(
      ins => gate6_outs,
      ins_valid => gate6_outs_valid,
      ins_ready => gate6_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork47_outs_0,
      outs(1) => fork47_outs_1,
      outs_valid(0) => fork47_outs_0_valid,
      outs_valid(1) => fork47_outs_1_valid,
      outs_ready(0) => fork47_outs_0_ready,
      outs_ready(1) => fork47_outs_1_ready
    );

  cmpi9 : entity work.handshake_cmpi_0(arch) generic map(32)
    port map(
      lhs => fork47_outs_1,
      lhs_valid => fork47_outs_1_valid,
      lhs_ready => fork47_outs_1_ready,
      rhs => extsi25_outs,
      rhs_valid => extsi25_outs_valid,
      rhs_ready => extsi25_outs_ready,
      clk => clk,
      rst => rst,
      result => cmpi9_result,
      result_valid => cmpi9_result_valid,
      result_ready => cmpi9_result_ready
    );

  fork48 : entity work.handshake_fork(arch) generic map(2, 1)
    port map(
      ins => cmpi9_result,
      ins_valid => cmpi9_result_valid,
      ins_ready => cmpi9_result_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork48_outs_0,
      outs(1) => fork48_outs_1,
      outs_valid(0) => fork48_outs_0_valid,
      outs_valid(1) => fork48_outs_1_valid,
      outs_ready(0) => fork48_outs_0_ready,
      outs_ready(1) => fork48_outs_1_ready
    );

  cmpi10 : entity work.handshake_cmpi_0(arch) generic map(32)
    port map(
      lhs => fork47_outs_0,
      lhs_valid => fork47_outs_0_valid,
      lhs_ready => fork47_outs_0_ready,
      rhs => fork11_outs_0,
      rhs_valid => fork11_outs_0_valid,
      rhs_ready => fork11_outs_0_ready,
      clk => clk,
      rst => rst,
      result => cmpi10_result,
      result_valid => cmpi10_result_valid,
      result_ready => cmpi10_result_ready
    );

  fork49 : entity work.handshake_fork(arch) generic map(2, 1)
    port map(
      ins => cmpi10_result,
      ins_valid => cmpi10_result_valid,
      ins_ready => cmpi10_result_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork49_outs_0,
      outs(1) => fork49_outs_1,
      outs_valid(0) => fork49_outs_0_valid,
      outs_valid(1) => fork49_outs_1_valid,
      outs_ready(0) => fork49_outs_0_ready,
      outs_ready(1) => fork49_outs_1_ready
    );

  cond_br95 : entity work.cond_br_dataless(arch)
    port map(
      condition => fork48_outs_1,
      condition_valid => fork48_outs_1_valid,
      condition_ready => fork48_outs_1_ready,
      data_valid => fork5_outs_1_valid,
      data_ready => fork5_outs_1_ready,
      clk => clk,
      rst => rst,
      trueOut_valid => cond_br95_trueOut_valid,
      trueOut_ready => cond_br95_trueOut_ready,
      falseOut_valid => cond_br95_falseOut_valid,
      falseOut_ready => cond_br95_falseOut_ready
    );

  sink35 : entity work.sink_dataless(arch)
    port map(
      ins_valid => cond_br95_trueOut_valid,
      ins_ready => cond_br95_trueOut_ready,
      clk => clk,
      rst => rst
    );

  cond_br96 : entity work.cond_br_dataless(arch)
    port map(
      condition => fork49_outs_1,
      condition_valid => fork49_outs_1_valid,
      condition_ready => fork49_outs_1_ready,
      data_valid => fork5_outs_0_valid,
      data_ready => fork5_outs_0_ready,
      clk => clk,
      rst => rst,
      trueOut_valid => cond_br96_trueOut_valid,
      trueOut_ready => cond_br96_trueOut_ready,
      falseOut_valid => cond_br96_falseOut_valid,
      falseOut_ready => cond_br96_falseOut_ready
    );

  sink36 : entity work.sink_dataless(arch)
    port map(
      ins_valid => cond_br96_trueOut_valid,
      ins_ready => cond_br96_trueOut_ready,
      clk => clk,
      rst => rst
    );

  source13 : entity work.source(arch)
    port map(
      clk => clk,
      rst => rst,
      outs_valid => source13_outs_valid,
      outs_ready => source13_outs_ready
    );

  mux91 : entity work.mux_dataless(arch) generic map(2, 1)
    port map(
      index => fork48_outs_0,
      index_valid => fork48_outs_0_valid,
      index_ready => fork48_outs_0_ready,
      ins_valid(0) => cond_br95_falseOut_valid,
      ins_valid(1) => source13_outs_valid,
      ins_ready(0) => cond_br95_falseOut_ready,
      ins_ready(1) => source13_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => mux91_outs_valid,
      outs_ready => mux91_outs_ready
    );

  source14 : entity work.source(arch)
    port map(
      clk => clk,
      rst => rst,
      outs_valid => source14_outs_valid,
      outs_ready => source14_outs_ready
    );

  mux92 : entity work.mux_dataless(arch) generic map(2, 1)
    port map(
      index => fork49_outs_0,
      index_valid => fork49_outs_0_valid,
      index_ready => fork49_outs_0_ready,
      ins_valid(0) => cond_br96_falseOut_valid,
      ins_valid(1) => source14_outs_valid,
      ins_ready(0) => cond_br96_falseOut_ready,
      ins_ready(1) => source14_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => mux92_outs_valid,
      outs_ready => mux92_outs_ready
    );

  buffer50 : entity work.tehb_dataless(arch)
    port map(
      ins_valid => mux91_outs_valid,
      ins_ready => mux91_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer50_outs_valid,
      outs_ready => buffer50_outs_ready
    );

  buffer51 : entity work.tehb_dataless(arch)
    port map(
      ins_valid => mux92_outs_valid,
      ins_ready => mux92_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer51_outs_valid,
      outs_ready => buffer51_outs_ready
    );

  join3 : entity work.join_handshake(arch) generic map(2)
    port map(
      ins_valid(0) => buffer50_outs_valid,
      ins_valid(1) => buffer51_outs_valid,
      ins_ready(0) => buffer50_outs_ready,
      ins_ready(1) => buffer51_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => join3_outs_valid,
      outs_ready => join3_outs_ready
    );

  buffer52 : entity work.oehb_dataless(arch)
    port map(
      ins_valid => join3_outs_valid,
      ins_ready => join3_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer52_outs_valid,
      outs_ready => buffer52_outs_ready
    );

  gate7 : entity work.gate(arch) generic map(2, 32)
    port map(
      ins(0) => buffer148_outs,
      ins_valid(0) => buffer148_outs_valid,
      ins_valid(1) => buffer52_outs_valid,
      ins_ready(0) => buffer148_outs_ready,
      ins_ready(1) => buffer52_outs_ready,
      clk => clk,
      rst => rst,
      outs => gate7_outs,
      outs_valid => gate7_outs_valid,
      outs_ready => gate7_outs_ready
    );

  buffer148 : entity work.tfifo(arch) generic map(1, 32)
    port map(
      ins => fork15_outs_4,
      ins_valid => fork15_outs_4_valid,
      ins_ready => fork15_outs_4_ready,
      clk => clk,
      rst => rst,
      outs => buffer148_outs,
      outs_valid => buffer148_outs_valid,
      outs_ready => buffer148_outs_ready
    );

  trunci3 : entity work.trunci(arch) generic map(32, 7)
    port map(
      ins => gate7_outs,
      ins_valid => gate7_outs_valid,
      ins_ready => gate7_outs_ready,
      clk => clk,
      rst => rst,
      outs => trunci3_outs,
      outs_valid => trunci3_outs_valid,
      outs_ready => trunci3_outs_ready
    );

  store0 : entity work.store(arch) generic map(32, 7)
    port map(
      addrIn => trunci3_outs,
      addrIn_valid => trunci3_outs_valid,
      addrIn_ready => trunci3_outs_ready,
      dataIn => addi7_result,
      dataIn_valid => addi7_result_valid,
      dataIn_ready => addi7_result_ready,
      doneFromMem_valid => mem_controller0_stDone_0_valid,
      doneFromMem_ready => mem_controller0_stDone_0_ready,
      clk => clk,
      rst => rst,
      addrOut => store0_addrOut,
      addrOut_valid => store0_addrOut_valid,
      addrOut_ready => store0_addrOut_ready,
      dataToMem => store0_dataToMem,
      dataToMem_valid => store0_dataToMem_valid,
      dataToMem_ready => store0_dataToMem_ready,
      doneOut_valid => store0_doneOut_valid,
      doneOut_ready => store0_doneOut_ready
    );

  addi4 : entity work.addi(arch) generic map(9)
    port map(
      lhs => extsi26_outs,
      lhs_valid => extsi26_outs_valid,
      lhs_ready => extsi26_outs_ready,
      rhs => extsi29_outs,
      rhs_valid => extsi29_outs_valid,
      rhs_ready => extsi29_outs_ready,
      clk => clk,
      rst => rst,
      result => addi4_result,
      result_valid => addi4_result_valid,
      result_ready => addi4_result_ready
    );

  buffer54 : entity work.oehb(arch) generic map(9)
    port map(
      ins => addi4_result,
      ins_valid => addi4_result_valid,
      ins_ready => addi4_result_ready,
      clk => clk,
      rst => rst,
      outs => buffer54_outs,
      outs_valid => buffer54_outs_valid,
      outs_ready => buffer54_outs_ready
    );

  fork50 : entity work.handshake_fork(arch) generic map(2, 9)
    port map(
      ins => buffer54_outs,
      ins_valid => buffer54_outs_valid,
      ins_ready => buffer54_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork50_outs_0,
      outs(1) => fork50_outs_1,
      outs_valid(0) => fork50_outs_0_valid,
      outs_valid(1) => fork50_outs_1_valid,
      outs_ready(0) => fork50_outs_0_ready,
      outs_ready(1) => fork50_outs_1_ready
    );

  trunci4 : entity work.trunci(arch) generic map(9, 8)
    port map(
      ins => fork50_outs_0,
      ins_valid => fork50_outs_0_valid,
      ins_ready => fork50_outs_0_ready,
      clk => clk,
      rst => rst,
      outs => trunci4_outs,
      outs_valid => trunci4_outs_valid,
      outs_ready => trunci4_outs_ready
    );

  cmpi0 : entity work.handshake_cmpi_1(arch) generic map(9)
    port map(
      lhs => fork50_outs_1,
      lhs_valid => fork50_outs_1_valid,
      lhs_ready => fork50_outs_1_ready,
      rhs => extsi31_outs,
      rhs_valid => extsi31_outs_valid,
      rhs_ready => extsi31_outs_ready,
      clk => clk,
      rst => rst,
      result => cmpi0_result,
      result_valid => cmpi0_result_valid,
      result_ready => cmpi0_result_ready
    );

  fork51 : entity work.handshake_fork(arch) generic map(34, 1)
    port map(
      ins => cmpi0_result,
      ins_valid => cmpi0_result_valid,
      ins_ready => cmpi0_result_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork51_outs_0,
      outs(1) => fork51_outs_1,
      outs(2) => fork51_outs_2,
      outs(3) => fork51_outs_3,
      outs(4) => fork51_outs_4,
      outs(5) => fork51_outs_5,
      outs(6) => fork51_outs_6,
      outs(7) => fork51_outs_7,
      outs(8) => fork51_outs_8,
      outs(9) => fork51_outs_9,
      outs(10) => fork51_outs_10,
      outs(11) => fork51_outs_11,
      outs(12) => fork51_outs_12,
      outs(13) => fork51_outs_13,
      outs(14) => fork51_outs_14,
      outs(15) => fork51_outs_15,
      outs(16) => fork51_outs_16,
      outs(17) => fork51_outs_17,
      outs(18) => fork51_outs_18,
      outs(19) => fork51_outs_19,
      outs(20) => fork51_outs_20,
      outs(21) => fork51_outs_21,
      outs(22) => fork51_outs_22,
      outs(23) => fork51_outs_23,
      outs(24) => fork51_outs_24,
      outs(25) => fork51_outs_25,
      outs(26) => fork51_outs_26,
      outs(27) => fork51_outs_27,
      outs(28) => fork51_outs_28,
      outs(29) => fork51_outs_29,
      outs(30) => fork51_outs_30,
      outs(31) => fork51_outs_31,
      outs(32) => fork51_outs_32,
      outs(33) => fork51_outs_33,
      outs_valid(0) => fork51_outs_0_valid,
      outs_valid(1) => fork51_outs_1_valid,
      outs_valid(2) => fork51_outs_2_valid,
      outs_valid(3) => fork51_outs_3_valid,
      outs_valid(4) => fork51_outs_4_valid,
      outs_valid(5) => fork51_outs_5_valid,
      outs_valid(6) => fork51_outs_6_valid,
      outs_valid(7) => fork51_outs_7_valid,
      outs_valid(8) => fork51_outs_8_valid,
      outs_valid(9) => fork51_outs_9_valid,
      outs_valid(10) => fork51_outs_10_valid,
      outs_valid(11) => fork51_outs_11_valid,
      outs_valid(12) => fork51_outs_12_valid,
      outs_valid(13) => fork51_outs_13_valid,
      outs_valid(14) => fork51_outs_14_valid,
      outs_valid(15) => fork51_outs_15_valid,
      outs_valid(16) => fork51_outs_16_valid,
      outs_valid(17) => fork51_outs_17_valid,
      outs_valid(18) => fork51_outs_18_valid,
      outs_valid(19) => fork51_outs_19_valid,
      outs_valid(20) => fork51_outs_20_valid,
      outs_valid(21) => fork51_outs_21_valid,
      outs_valid(22) => fork51_outs_22_valid,
      outs_valid(23) => fork51_outs_23_valid,
      outs_valid(24) => fork51_outs_24_valid,
      outs_valid(25) => fork51_outs_25_valid,
      outs_valid(26) => fork51_outs_26_valid,
      outs_valid(27) => fork51_outs_27_valid,
      outs_valid(28) => fork51_outs_28_valid,
      outs_valid(29) => fork51_outs_29_valid,
      outs_valid(30) => fork51_outs_30_valid,
      outs_valid(31) => fork51_outs_31_valid,
      outs_valid(32) => fork51_outs_32_valid,
      outs_valid(33) => fork51_outs_33_valid,
      outs_ready(0) => fork51_outs_0_ready,
      outs_ready(1) => fork51_outs_1_ready,
      outs_ready(2) => fork51_outs_2_ready,
      outs_ready(3) => fork51_outs_3_ready,
      outs_ready(4) => fork51_outs_4_ready,
      outs_ready(5) => fork51_outs_5_ready,
      outs_ready(6) => fork51_outs_6_ready,
      outs_ready(7) => fork51_outs_7_ready,
      outs_ready(8) => fork51_outs_8_ready,
      outs_ready(9) => fork51_outs_9_ready,
      outs_ready(10) => fork51_outs_10_ready,
      outs_ready(11) => fork51_outs_11_ready,
      outs_ready(12) => fork51_outs_12_ready,
      outs_ready(13) => fork51_outs_13_ready,
      outs_ready(14) => fork51_outs_14_ready,
      outs_ready(15) => fork51_outs_15_ready,
      outs_ready(16) => fork51_outs_16_ready,
      outs_ready(17) => fork51_outs_17_ready,
      outs_ready(18) => fork51_outs_18_ready,
      outs_ready(19) => fork51_outs_19_ready,
      outs_ready(20) => fork51_outs_20_ready,
      outs_ready(21) => fork51_outs_21_ready,
      outs_ready(22) => fork51_outs_22_ready,
      outs_ready(23) => fork51_outs_23_ready,
      outs_ready(24) => fork51_outs_24_ready,
      outs_ready(25) => fork51_outs_25_ready,
      outs_ready(26) => fork51_outs_26_ready,
      outs_ready(27) => fork51_outs_27_ready,
      outs_ready(28) => fork51_outs_28_ready,
      outs_ready(29) => fork51_outs_29_ready,
      outs_ready(30) => fork51_outs_30_ready,
      outs_ready(31) => fork51_outs_31_ready,
      outs_ready(32) => fork51_outs_32_ready,
      outs_ready(33) => fork51_outs_33_ready
    );

  cond_br3 : entity work.cond_br(arch) generic map(8)
    port map(
      condition => fork51_outs_0,
      condition_valid => fork51_outs_0_valid,
      condition_ready => fork51_outs_0_ready,
      data => trunci4_outs,
      data_valid => trunci4_outs_valid,
      data_ready => trunci4_outs_ready,
      clk => clk,
      rst => rst,
      trueOut => cond_br3_trueOut,
      trueOut_valid => cond_br3_trueOut_valid,
      trueOut_ready => cond_br3_trueOut_ready,
      falseOut => cond_br3_falseOut,
      falseOut_valid => cond_br3_falseOut_valid,
      falseOut_ready => cond_br3_falseOut_ready
    );

  sink37 : entity work.sink(arch) generic map(8)
    port map(
      ins => cond_br3_falseOut,
      ins_valid => cond_br3_falseOut_valid,
      ins_ready => cond_br3_falseOut_ready,
      clk => clk,
      rst => rst
    );

  buffer34 : entity work.oehb(arch) generic map(3)
    port map(
      ins => mux2_outs,
      ins_valid => mux2_outs_valid,
      ins_ready => mux2_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer34_outs,
      outs_valid => buffer34_outs_valid,
      outs_ready => buffer34_outs_ready
    );

  buffer35 : entity work.tehb(arch) generic map(3)
    port map(
      ins => buffer34_outs,
      ins_valid => buffer34_outs_valid,
      ins_ready => buffer34_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer35_outs,
      outs_valid => buffer35_outs_valid,
      outs_ready => buffer35_outs_ready
    );

  cond_br4 : entity work.cond_br(arch) generic map(3)
    port map(
      condition => fork51_outs_5,
      condition_valid => fork51_outs_5_valid,
      condition_ready => fork51_outs_5_ready,
      data => buffer35_outs,
      data_valid => buffer35_outs_valid,
      data_ready => buffer35_outs_ready,
      clk => clk,
      rst => rst,
      trueOut => cond_br4_trueOut,
      trueOut_valid => cond_br4_trueOut_valid,
      trueOut_ready => cond_br4_trueOut_ready,
      falseOut => cond_br4_falseOut,
      falseOut_valid => cond_br4_falseOut_valid,
      falseOut_ready => cond_br4_falseOut_ready
    );

  cond_br5 : entity work.cond_br_dataless(arch)
    port map(
      condition => fork51_outs_32,
      condition_valid => fork51_outs_32_valid,
      condition_ready => fork51_outs_32_ready,
      data_valid => fork17_outs_1_valid,
      data_ready => fork17_outs_1_ready,
      clk => clk,
      rst => rst,
      trueOut_valid => cond_br5_trueOut_valid,
      trueOut_ready => cond_br5_trueOut_ready,
      falseOut_valid => cond_br5_falseOut_valid,
      falseOut_ready => cond_br5_falseOut_ready
    );

  cond_br6 : entity work.cond_br(arch) generic map(2)
    port map(
      condition => fork51_outs_33,
      condition_valid => fork51_outs_33_valid,
      condition_ready => fork51_outs_33_ready,
      data => fork18_outs_2,
      data_valid => fork18_outs_2_valid,
      data_ready => fork18_outs_2_ready,
      clk => clk,
      rst => rst,
      trueOut => cond_br6_trueOut,
      trueOut_valid => cond_br6_trueOut_valid,
      trueOut_ready => cond_br6_trueOut_ready,
      falseOut => cond_br6_falseOut,
      falseOut_valid => cond_br6_falseOut_valid,
      falseOut_ready => cond_br6_falseOut_ready
    );

  sink38 : entity work.sink(arch) generic map(2)
    port map(
      ins => cond_br6_trueOut,
      ins_valid => cond_br6_trueOut_valid,
      ins_ready => cond_br6_trueOut_ready,
      clk => clk,
      rst => rst
    );

  extsi19 : entity work.extsi(arch) generic map(2, 8)
    port map(
      ins => cond_br6_falseOut,
      ins_valid => cond_br6_falseOut_valid,
      ins_ready => cond_br6_falseOut_ready,
      clk => clk,
      rst => rst,
      outs => extsi19_outs,
      outs_valid => extsi19_outs_valid,
      outs_ready => extsi19_outs_ready
    );

  cond_br234 : entity work.cond_br(arch) generic map(9)
    port map(
      condition => fork94_outs_3,
      condition_valid => fork94_outs_3_valid,
      condition_ready => fork94_outs_3_ready,
      data => fork57_outs_0,
      data_valid => fork57_outs_0_valid,
      data_ready => fork57_outs_0_ready,
      clk => clk,
      rst => rst,
      trueOut => cond_br234_trueOut,
      trueOut_valid => cond_br234_trueOut_valid,
      trueOut_ready => cond_br234_trueOut_ready,
      falseOut => cond_br234_falseOut,
      falseOut_valid => cond_br234_falseOut_valid,
      falseOut_ready => cond_br234_falseOut_ready
    );

  sink39 : entity work.sink(arch) generic map(9)
    port map(
      ins => cond_br234_falseOut,
      ins_valid => cond_br234_falseOut_valid,
      ins_ready => cond_br234_falseOut_ready,
      clk => clk,
      rst => rst
    );

  cond_br235 : entity work.cond_br(arch) generic map(32)
    port map(
      condition => fork94_outs_27,
      condition_valid => fork94_outs_27_valid,
      condition_ready => fork94_outs_27_ready,
      data => fork70_outs_1,
      data_valid => fork70_outs_1_valid,
      data_ready => fork70_outs_1_ready,
      clk => clk,
      rst => rst,
      trueOut => cond_br235_trueOut,
      trueOut_valid => cond_br235_trueOut_valid,
      trueOut_ready => cond_br235_trueOut_ready,
      falseOut => cond_br235_falseOut,
      falseOut_valid => cond_br235_falseOut_valid,
      falseOut_ready => cond_br235_falseOut_ready
    );

  sink40 : entity work.sink(arch) generic map(32)
    port map(
      ins => cond_br235_falseOut,
      ins_valid => cond_br235_falseOut_valid,
      ins_ready => cond_br235_falseOut_ready,
      clk => clk,
      rst => rst
    );

  cond_br236 : entity work.cond_br_dataless(arch)
    port map(
      condition => buffer160_outs,
      condition_valid => buffer160_outs_valid,
      condition_ready => buffer160_outs_ready,
      data_valid => fork62_outs_1_valid,
      data_ready => fork62_outs_1_ready,
      clk => clk,
      rst => rst,
      trueOut_valid => cond_br236_trueOut_valid,
      trueOut_ready => cond_br236_trueOut_ready,
      falseOut_valid => cond_br236_falseOut_valid,
      falseOut_ready => cond_br236_falseOut_ready
    );

  buffer160 : entity work.tfifo(arch) generic map(1, 1)
    port map(
      ins => fork94_outs_26,
      ins_valid => fork94_outs_26_valid,
      ins_ready => fork94_outs_26_ready,
      clk => clk,
      rst => rst,
      outs => buffer160_outs,
      outs_valid => buffer160_outs_valid,
      outs_ready => buffer160_outs_ready
    );

  sink41 : entity work.sink_dataless(arch)
    port map(
      ins_valid => cond_br236_falseOut_valid,
      ins_ready => cond_br236_falseOut_ready,
      clk => clk,
      rst => rst
    );

  cond_br237 : entity work.cond_br_dataless(arch)
    port map(
      condition => fork94_outs_25,
      condition_valid => fork94_outs_25_valid,
      condition_ready => fork94_outs_25_ready,
      data_valid => fork61_outs_1_valid,
      data_ready => fork61_outs_1_ready,
      clk => clk,
      rst => rst,
      trueOut_valid => cond_br237_trueOut_valid,
      trueOut_ready => cond_br237_trueOut_ready,
      falseOut_valid => cond_br237_falseOut_valid,
      falseOut_ready => cond_br237_falseOut_ready
    );

  sink42 : entity work.sink_dataless(arch)
    port map(
      ins_valid => cond_br237_falseOut_valid,
      ins_ready => cond_br237_falseOut_ready,
      clk => clk,
      rst => rst
    );

  cond_br238 : entity work.cond_br_dataless(arch)
    port map(
      condition => fork94_outs_24,
      condition_valid => fork94_outs_24_valid,
      condition_ready => fork94_outs_24_ready,
      data_valid => fork64_outs_1_valid,
      data_ready => fork64_outs_1_ready,
      clk => clk,
      rst => rst,
      trueOut_valid => cond_br238_trueOut_valid,
      trueOut_ready => cond_br238_trueOut_ready,
      falseOut_valid => cond_br238_falseOut_valid,
      falseOut_ready => cond_br238_falseOut_ready
    );

  sink43 : entity work.sink_dataless(arch)
    port map(
      ins_valid => cond_br238_falseOut_valid,
      ins_ready => cond_br238_falseOut_ready,
      clk => clk,
      rst => rst
    );

  cond_br239 : entity work.cond_br(arch) generic map(32)
    port map(
      condition => fork94_outs_23,
      condition_valid => fork94_outs_23_valid,
      condition_ready => fork94_outs_23_ready,
      data => fork59_outs_1,
      data_valid => fork59_outs_1_valid,
      data_ready => fork59_outs_1_ready,
      clk => clk,
      rst => rst,
      trueOut => cond_br239_trueOut,
      trueOut_valid => cond_br239_trueOut_valid,
      trueOut_ready => cond_br239_trueOut_ready,
      falseOut => cond_br239_falseOut,
      falseOut_valid => cond_br239_falseOut_valid,
      falseOut_ready => cond_br239_falseOut_ready
    );

  sink44 : entity work.sink(arch) generic map(32)
    port map(
      ins => cond_br239_falseOut,
      ins_valid => cond_br239_falseOut_valid,
      ins_ready => cond_br239_falseOut_ready,
      clk => clk,
      rst => rst
    );

  cond_br240 : entity work.cond_br_dataless(arch)
    port map(
      condition => fork94_outs_22,
      condition_valid => fork94_outs_22_valid,
      condition_ready => fork94_outs_22_ready,
      data_valid => fork65_outs_1_valid,
      data_ready => fork65_outs_1_ready,
      clk => clk,
      rst => rst,
      trueOut_valid => cond_br240_trueOut_valid,
      trueOut_ready => cond_br240_trueOut_ready,
      falseOut_valid => cond_br240_falseOut_valid,
      falseOut_ready => cond_br240_falseOut_ready
    );

  sink45 : entity work.sink_dataless(arch)
    port map(
      ins_valid => cond_br240_falseOut_valid,
      ins_ready => cond_br240_falseOut_ready,
      clk => clk,
      rst => rst
    );

  cond_br241 : entity work.cond_br_dataless(arch)
    port map(
      condition => fork94_outs_21,
      condition_valid => fork94_outs_21_valid,
      condition_ready => fork94_outs_21_ready,
      data_valid => fork66_outs_1_valid,
      data_ready => fork66_outs_1_ready,
      clk => clk,
      rst => rst,
      trueOut_valid => cond_br241_trueOut_valid,
      trueOut_ready => cond_br241_trueOut_ready,
      falseOut_valid => cond_br241_falseOut_valid,
      falseOut_ready => cond_br241_falseOut_ready
    );

  sink46 : entity work.sink_dataless(arch)
    port map(
      ins_valid => cond_br241_falseOut_valid,
      ins_ready => cond_br241_falseOut_ready,
      clk => clk,
      rst => rst
    );

  cond_br242 : entity work.cond_br(arch) generic map(8)
    port map(
      condition => fork94_outs_2,
      condition_valid => fork94_outs_2_valid,
      condition_ready => fork94_outs_2_ready,
      data => fork58_outs_0,
      data_valid => fork58_outs_0_valid,
      data_ready => fork58_outs_0_ready,
      clk => clk,
      rst => rst,
      trueOut => cond_br242_trueOut,
      trueOut_valid => cond_br242_trueOut_valid,
      trueOut_ready => cond_br242_trueOut_ready,
      falseOut => cond_br242_falseOut,
      falseOut_valid => cond_br242_falseOut_valid,
      falseOut_ready => cond_br242_falseOut_ready
    );

  sink47 : entity work.sink(arch) generic map(8)
    port map(
      ins => cond_br242_falseOut,
      ins_valid => cond_br242_falseOut_valid,
      ins_ready => cond_br242_falseOut_ready,
      clk => clk,
      rst => rst
    );

  cond_br243 : entity work.cond_br_dataless(arch)
    port map(
      condition => fork94_outs_20,
      condition_valid => fork94_outs_20_valid,
      condition_ready => fork94_outs_20_ready,
      data_valid => fork71_outs_1_valid,
      data_ready => fork71_outs_1_ready,
      clk => clk,
      rst => rst,
      trueOut_valid => cond_br243_trueOut_valid,
      trueOut_ready => cond_br243_trueOut_ready,
      falseOut_valid => cond_br243_falseOut_valid,
      falseOut_ready => cond_br243_falseOut_ready
    );

  sink48 : entity work.sink_dataless(arch)
    port map(
      ins_valid => cond_br243_falseOut_valid,
      ins_ready => cond_br243_falseOut_ready,
      clk => clk,
      rst => rst
    );

  cond_br244 : entity work.cond_br(arch) generic map(32)
    port map(
      condition => fork94_outs_19,
      condition_valid => fork94_outs_19_valid,
      condition_ready => fork94_outs_19_ready,
      data => init135_outs,
      data_valid => init135_outs_valid,
      data_ready => init135_outs_ready,
      clk => clk,
      rst => rst,
      trueOut => cond_br244_trueOut,
      trueOut_valid => cond_br244_trueOut_valid,
      trueOut_ready => cond_br244_trueOut_ready,
      falseOut => cond_br244_falseOut,
      falseOut_valid => cond_br244_falseOut_valid,
      falseOut_ready => cond_br244_falseOut_ready
    );

  sink49 : entity work.sink(arch) generic map(32)
    port map(
      ins => cond_br244_trueOut,
      ins_valid => cond_br244_trueOut_valid,
      ins_ready => cond_br244_trueOut_ready,
      clk => clk,
      rst => rst
    );

  cond_br245 : entity work.cond_br_dataless(arch)
    port map(
      condition => fork94_outs_18,
      condition_valid => fork94_outs_18_valid,
      condition_ready => fork94_outs_18_ready,
      data_valid => fork72_outs_1_valid,
      data_ready => fork72_outs_1_ready,
      clk => clk,
      rst => rst,
      trueOut_valid => cond_br245_trueOut_valid,
      trueOut_ready => cond_br245_trueOut_ready,
      falseOut_valid => cond_br245_falseOut_valid,
      falseOut_ready => cond_br245_falseOut_ready
    );

  sink50 : entity work.sink_dataless(arch)
    port map(
      ins_valid => cond_br245_falseOut_valid,
      ins_ready => cond_br245_falseOut_ready,
      clk => clk,
      rst => rst
    );

  cond_br246 : entity work.cond_br(arch) generic map(8)
    port map(
      condition => fork94_outs_5,
      condition_valid => fork94_outs_5_valid,
      condition_ready => fork94_outs_5_ready,
      data => fork91_outs_0,
      data_valid => fork91_outs_0_valid,
      data_ready => fork91_outs_0_ready,
      clk => clk,
      rst => rst,
      trueOut => cond_br246_trueOut,
      trueOut_valid => cond_br246_trueOut_valid,
      trueOut_ready => cond_br246_trueOut_ready,
      falseOut => cond_br246_falseOut,
      falseOut_valid => cond_br246_falseOut_valid,
      falseOut_ready => cond_br246_falseOut_ready
    );

  sink51 : entity work.sink(arch) generic map(8)
    port map(
      ins => cond_br246_trueOut,
      ins_valid => cond_br246_trueOut_valid,
      ins_ready => cond_br246_trueOut_ready,
      clk => clk,
      rst => rst
    );

  cond_br247 : entity work.cond_br_dataless(arch)
    port map(
      condition => buffer174_outs,
      condition_valid => buffer174_outs_valid,
      condition_ready => buffer174_outs_ready,
      data_valid => fork67_outs_1_valid,
      data_ready => fork67_outs_1_ready,
      clk => clk,
      rst => rst,
      trueOut_valid => cond_br247_trueOut_valid,
      trueOut_ready => cond_br247_trueOut_ready,
      falseOut_valid => cond_br247_falseOut_valid,
      falseOut_ready => cond_br247_falseOut_ready
    );

  buffer174 : entity work.tfifo(arch) generic map(1, 1)
    port map(
      ins => fork94_outs_17,
      ins_valid => fork94_outs_17_valid,
      ins_ready => fork94_outs_17_ready,
      clk => clk,
      rst => rst,
      outs => buffer174_outs,
      outs_valid => buffer174_outs_valid,
      outs_ready => buffer174_outs_ready
    );

  sink52 : entity work.sink_dataless(arch)
    port map(
      ins_valid => cond_br247_falseOut_valid,
      ins_ready => cond_br247_falseOut_ready,
      clk => clk,
      rst => rst
    );

  cond_br248 : entity work.cond_br_dataless(arch)
    port map(
      condition => buffer175_outs,
      condition_valid => buffer175_outs_valid,
      condition_ready => buffer175_outs_ready,
      data_valid => fork60_outs_1_valid,
      data_ready => fork60_outs_1_ready,
      clk => clk,
      rst => rst,
      trueOut_valid => cond_br248_trueOut_valid,
      trueOut_ready => cond_br248_trueOut_ready,
      falseOut_valid => cond_br248_falseOut_valid,
      falseOut_ready => cond_br248_falseOut_ready
    );

  buffer175 : entity work.tfifo(arch) generic map(1, 1)
    port map(
      ins => fork94_outs_16,
      ins_valid => fork94_outs_16_valid,
      ins_ready => fork94_outs_16_ready,
      clk => clk,
      rst => rst,
      outs => buffer175_outs,
      outs_valid => buffer175_outs_valid,
      outs_ready => buffer175_outs_ready
    );

  sink53 : entity work.sink_dataless(arch)
    port map(
      ins_valid => cond_br248_falseOut_valid,
      ins_ready => cond_br248_falseOut_ready,
      clk => clk,
      rst => rst
    );

  cond_br249 : entity work.cond_br(arch) generic map(32)
    port map(
      condition => fork94_outs_15,
      condition_valid => fork94_outs_15_valid,
      condition_ready => fork94_outs_15_ready,
      data => init132_outs,
      data_valid => init132_outs_valid,
      data_ready => init132_outs_ready,
      clk => clk,
      rst => rst,
      trueOut => cond_br249_trueOut,
      trueOut_valid => cond_br249_trueOut_valid,
      trueOut_ready => cond_br249_trueOut_ready,
      falseOut => cond_br249_falseOut,
      falseOut_valid => cond_br249_falseOut_valid,
      falseOut_ready => cond_br249_falseOut_ready
    );

  sink54 : entity work.sink(arch) generic map(32)
    port map(
      ins => cond_br249_trueOut,
      ins_valid => cond_br249_trueOut_valid,
      ins_ready => cond_br249_trueOut_ready,
      clk => clk,
      rst => rst
    );

  cond_br250 : entity work.cond_br_dataless(arch)
    port map(
      condition => buffer177_outs,
      condition_valid => buffer177_outs_valid,
      condition_ready => buffer177_outs_ready,
      data_valid => fork54_outs_1_valid,
      data_ready => fork54_outs_1_ready,
      clk => clk,
      rst => rst,
      trueOut_valid => cond_br250_trueOut_valid,
      trueOut_ready => cond_br250_trueOut_ready,
      falseOut_valid => cond_br250_falseOut_valid,
      falseOut_ready => cond_br250_falseOut_ready
    );

  buffer177 : entity work.tfifo(arch) generic map(1, 1)
    port map(
      ins => fork94_outs_14,
      ins_valid => fork94_outs_14_valid,
      ins_ready => fork94_outs_14_ready,
      clk => clk,
      rst => rst,
      outs => buffer177_outs,
      outs_valid => buffer177_outs_valid,
      outs_ready => buffer177_outs_ready
    );

  sink55 : entity work.sink_dataless(arch)
    port map(
      ins_valid => cond_br250_falseOut_valid,
      ins_ready => cond_br250_falseOut_ready,
      clk => clk,
      rst => rst
    );

  cond_br251 : entity work.cond_br(arch) generic map(32)
    port map(
      condition => fork94_outs_13,
      condition_valid => fork94_outs_13_valid,
      condition_ready => fork94_outs_13_ready,
      data => buffer179_outs,
      data_valid => buffer179_outs_valid,
      data_ready => buffer179_outs_ready,
      clk => clk,
      rst => rst,
      trueOut => cond_br251_trueOut,
      trueOut_valid => cond_br251_trueOut_valid,
      trueOut_ready => cond_br251_trueOut_ready,
      falseOut => cond_br251_falseOut,
      falseOut_valid => cond_br251_falseOut_valid,
      falseOut_ready => cond_br251_falseOut_ready
    );

  buffer179 : entity work.tfifo(arch) generic map(1, 32)
    port map(
      ins => fork55_outs_1,
      ins_valid => fork55_outs_1_valid,
      ins_ready => fork55_outs_1_ready,
      clk => clk,
      rst => rst,
      outs => buffer179_outs,
      outs_valid => buffer179_outs_valid,
      outs_ready => buffer179_outs_ready
    );

  sink56 : entity work.sink(arch) generic map(32)
    port map(
      ins => cond_br251_falseOut,
      ins_valid => cond_br251_falseOut_valid,
      ins_ready => cond_br251_falseOut_ready,
      clk => clk,
      rst => rst
    );

  cond_br252 : entity work.cond_br(arch) generic map(8)
    port map(
      condition => buffer180_outs,
      condition_valid => buffer180_outs_valid,
      condition_ready => buffer180_outs_ready,
      data => fork53_outs_0,
      data_valid => fork53_outs_0_valid,
      data_ready => fork53_outs_0_ready,
      clk => clk,
      rst => rst,
      trueOut => cond_br252_trueOut,
      trueOut_valid => cond_br252_trueOut_valid,
      trueOut_ready => cond_br252_trueOut_ready,
      falseOut => cond_br252_falseOut,
      falseOut_valid => cond_br252_falseOut_valid,
      falseOut_ready => cond_br252_falseOut_ready
    );

  buffer180 : entity work.tfifo(arch) generic map(1, 1)
    port map(
      ins => fork94_outs_4,
      ins_valid => fork94_outs_4_valid,
      ins_ready => fork94_outs_4_ready,
      clk => clk,
      rst => rst,
      outs => buffer180_outs,
      outs_valid => buffer180_outs_valid,
      outs_ready => buffer180_outs_ready
    );

  sink57 : entity work.sink(arch) generic map(8)
    port map(
      ins => cond_br252_falseOut,
      ins_valid => cond_br252_falseOut_valid,
      ins_ready => cond_br252_falseOut_ready,
      clk => clk,
      rst => rst
    );

  cond_br253 : entity work.cond_br_dataless(arch)
    port map(
      condition => fork94_outs_12,
      condition_valid => fork94_outs_12_valid,
      condition_ready => fork94_outs_12_ready,
      data_valid => fork68_outs_1_valid,
      data_ready => fork68_outs_1_ready,
      clk => clk,
      rst => rst,
      trueOut_valid => cond_br253_trueOut_valid,
      trueOut_ready => cond_br253_trueOut_ready,
      falseOut_valid => cond_br253_falseOut_valid,
      falseOut_ready => cond_br253_falseOut_ready
    );

  sink58 : entity work.sink_dataless(arch)
    port map(
      ins_valid => cond_br253_falseOut_valid,
      ins_ready => cond_br253_falseOut_ready,
      clk => clk,
      rst => rst
    );

  cond_br254 : entity work.cond_br(arch) generic map(32)
    port map(
      condition => fork94_outs_11,
      condition_valid => fork94_outs_11_valid,
      condition_ready => fork94_outs_11_ready,
      data => buffer184_outs,
      data_valid => buffer184_outs_valid,
      data_ready => buffer184_outs_ready,
      clk => clk,
      rst => rst,
      trueOut => cond_br254_trueOut,
      trueOut_valid => cond_br254_trueOut_valid,
      trueOut_ready => cond_br254_trueOut_ready,
      falseOut => cond_br254_falseOut,
      falseOut_valid => cond_br254_falseOut_valid,
      falseOut_ready => cond_br254_falseOut_ready
    );

  buffer184 : entity work.tfifo(arch) generic map(1, 32)
    port map(
      ins => fork69_outs_1,
      ins_valid => fork69_outs_1_valid,
      ins_ready => fork69_outs_1_ready,
      clk => clk,
      rst => rst,
      outs => buffer184_outs,
      outs_valid => buffer184_outs_valid,
      outs_ready => buffer184_outs_ready
    );

  sink59 : entity work.sink(arch) generic map(32)
    port map(
      ins => cond_br254_falseOut,
      ins_valid => cond_br254_falseOut_valid,
      ins_ready => cond_br254_falseOut_ready,
      clk => clk,
      rst => rst
    );

  cond_br255 : entity work.cond_br_dataless(arch)
    port map(
      condition => buffer185_outs,
      condition_valid => buffer185_outs_valid,
      condition_ready => buffer185_outs_ready,
      data_valid => fork56_outs_1_valid,
      data_ready => fork56_outs_1_ready,
      clk => clk,
      rst => rst,
      trueOut_valid => cond_br255_trueOut_valid,
      trueOut_ready => cond_br255_trueOut_ready,
      falseOut_valid => cond_br255_falseOut_valid,
      falseOut_ready => cond_br255_falseOut_ready
    );

  buffer185 : entity work.tfifo(arch) generic map(1, 1)
    port map(
      ins => fork94_outs_10,
      ins_valid => fork94_outs_10_valid,
      ins_ready => fork94_outs_10_ready,
      clk => clk,
      rst => rst,
      outs => buffer185_outs,
      outs_valid => buffer185_outs_valid,
      outs_ready => buffer185_outs_ready
    );

  sink60 : entity work.sink_dataless(arch)
    port map(
      ins_valid => cond_br255_falseOut_valid,
      ins_ready => cond_br255_falseOut_ready,
      clk => clk,
      rst => rst
    );

  cond_br256 : entity work.cond_br(arch) generic map(32)
    port map(
      condition => buffer186_outs,
      condition_valid => buffer186_outs_valid,
      condition_ready => buffer186_outs_ready,
      data => buffer187_outs,
      data_valid => buffer187_outs_valid,
      data_ready => buffer187_outs_ready,
      clk => clk,
      rst => rst,
      trueOut => cond_br256_trueOut,
      trueOut_valid => cond_br256_trueOut_valid,
      trueOut_ready => cond_br256_trueOut_ready,
      falseOut => cond_br256_falseOut,
      falseOut_valid => cond_br256_falseOut_valid,
      falseOut_ready => cond_br256_falseOut_ready
    );

  buffer186 : entity work.tfifo(arch) generic map(1, 1)
    port map(
      ins => fork94_outs_9,
      ins_valid => fork94_outs_9_valid,
      ins_ready => fork94_outs_9_ready,
      clk => clk,
      rst => rst,
      outs => buffer186_outs,
      outs_valid => buffer186_outs_valid,
      outs_ready => buffer186_outs_ready
    );

  buffer187 : entity work.tfifo(arch) generic map(1, 32)
    port map(
      ins => fork63_outs_1,
      ins_valid => fork63_outs_1_valid,
      ins_ready => fork63_outs_1_ready,
      clk => clk,
      rst => rst,
      outs => buffer187_outs,
      outs_valid => buffer187_outs_valid,
      outs_ready => buffer187_outs_ready
    );

  sink61 : entity work.sink(arch) generic map(32)
    port map(
      ins => cond_br256_falseOut,
      ins_valid => cond_br256_falseOut_valid,
      ins_ready => cond_br256_falseOut_ready,
      clk => clk,
      rst => rst
    );

  cond_br257 : entity work.cond_br_dataless(arch)
    port map(
      condition => buffer188_outs,
      condition_valid => buffer188_outs_valid,
      condition_ready => buffer188_outs_ready,
      data_valid => fork92_outs_1_valid,
      data_ready => fork92_outs_1_ready,
      clk => clk,
      rst => rst,
      trueOut_valid => cond_br257_trueOut_valid,
      trueOut_ready => cond_br257_trueOut_ready,
      falseOut_valid => cond_br257_falseOut_valid,
      falseOut_ready => cond_br257_falseOut_ready
    );

  buffer188 : entity work.tfifo(arch) generic map(1, 1)
    port map(
      ins => fork94_outs_8,
      ins_valid => fork94_outs_8_valid,
      ins_ready => fork94_outs_8_ready,
      clk => clk,
      rst => rst,
      outs => buffer188_outs,
      outs_valid => buffer188_outs_valid,
      outs_ready => buffer188_outs_ready
    );

  sink62 : entity work.sink_dataless(arch)
    port map(
      ins_valid => cond_br257_trueOut_valid,
      ins_ready => cond_br257_trueOut_ready,
      clk => clk,
      rst => rst
    );

  cond_br258 : entity work.cond_br(arch) generic map(8)
    port map(
      condition => fork94_outs_6,
      condition_valid => fork94_outs_6_valid,
      condition_ready => fork94_outs_6_ready,
      data => fork80_outs_0,
      data_valid => fork80_outs_0_valid,
      data_ready => fork80_outs_0_ready,
      clk => clk,
      rst => rst,
      trueOut => cond_br258_trueOut,
      trueOut_valid => cond_br258_trueOut_valid,
      trueOut_ready => cond_br258_trueOut_ready,
      falseOut => cond_br258_falseOut,
      falseOut_valid => cond_br258_falseOut_valid,
      falseOut_ready => cond_br258_falseOut_ready
    );

  sink63 : entity work.sink(arch) generic map(8)
    port map(
      ins => cond_br258_trueOut,
      ins_valid => cond_br258_trueOut_valid,
      ins_ready => cond_br258_trueOut_ready,
      clk => clk,
      rst => rst
    );

  init92 : entity work.tehb_init(arch) generic map(1, 0)
    port map(
      ins => fork94_outs_7,
      ins_valid => fork94_outs_7_valid,
      ins_ready => fork94_outs_7_ready,
      clk => clk,
      rst => rst,
      outs => init92_outs,
      outs_valid => init92_outs_valid,
      outs_ready => init92_outs_ready
    );

  fork52 : entity work.handshake_fork(arch) generic map(20, 1)
    port map(
      ins => init92_outs,
      ins_valid => init92_outs_valid,
      ins_ready => init92_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork52_outs_0,
      outs(1) => fork52_outs_1,
      outs(2) => fork52_outs_2,
      outs(3) => fork52_outs_3,
      outs(4) => fork52_outs_4,
      outs(5) => fork52_outs_5,
      outs(6) => fork52_outs_6,
      outs(7) => fork52_outs_7,
      outs(8) => fork52_outs_8,
      outs(9) => fork52_outs_9,
      outs(10) => fork52_outs_10,
      outs(11) => fork52_outs_11,
      outs(12) => fork52_outs_12,
      outs(13) => fork52_outs_13,
      outs(14) => fork52_outs_14,
      outs(15) => fork52_outs_15,
      outs(16) => fork52_outs_16,
      outs(17) => fork52_outs_17,
      outs(18) => fork52_outs_18,
      outs(19) => fork52_outs_19,
      outs_valid(0) => fork52_outs_0_valid,
      outs_valid(1) => fork52_outs_1_valid,
      outs_valid(2) => fork52_outs_2_valid,
      outs_valid(3) => fork52_outs_3_valid,
      outs_valid(4) => fork52_outs_4_valid,
      outs_valid(5) => fork52_outs_5_valid,
      outs_valid(6) => fork52_outs_6_valid,
      outs_valid(7) => fork52_outs_7_valid,
      outs_valid(8) => fork52_outs_8_valid,
      outs_valid(9) => fork52_outs_9_valid,
      outs_valid(10) => fork52_outs_10_valid,
      outs_valid(11) => fork52_outs_11_valid,
      outs_valid(12) => fork52_outs_12_valid,
      outs_valid(13) => fork52_outs_13_valid,
      outs_valid(14) => fork52_outs_14_valid,
      outs_valid(15) => fork52_outs_15_valid,
      outs_valid(16) => fork52_outs_16_valid,
      outs_valid(17) => fork52_outs_17_valid,
      outs_valid(18) => fork52_outs_18_valid,
      outs_valid(19) => fork52_outs_19_valid,
      outs_ready(0) => fork52_outs_0_ready,
      outs_ready(1) => fork52_outs_1_ready,
      outs_ready(2) => fork52_outs_2_ready,
      outs_ready(3) => fork52_outs_3_ready,
      outs_ready(4) => fork52_outs_4_ready,
      outs_ready(5) => fork52_outs_5_ready,
      outs_ready(6) => fork52_outs_6_ready,
      outs_ready(7) => fork52_outs_7_ready,
      outs_ready(8) => fork52_outs_8_ready,
      outs_ready(9) => fork52_outs_9_ready,
      outs_ready(10) => fork52_outs_10_ready,
      outs_ready(11) => fork52_outs_11_ready,
      outs_ready(12) => fork52_outs_12_ready,
      outs_ready(13) => fork52_outs_13_ready,
      outs_ready(14) => fork52_outs_14_ready,
      outs_ready(15) => fork52_outs_15_ready,
      outs_ready(16) => fork52_outs_16_ready,
      outs_ready(17) => fork52_outs_17_ready,
      outs_ready(18) => fork52_outs_18_ready,
      outs_ready(19) => fork52_outs_19_ready
    );

  mux93 : entity work.mux(arch) generic map(2, 8, 1)
    port map(
      index => fork52_outs_2,
      index_valid => fork52_outs_2_valid,
      index_ready => fork52_outs_2_ready,
      ins(0) => cond_br230_falseOut,
      ins(1) => cond_br252_trueOut,
      ins_valid(0) => cond_br230_falseOut_valid,
      ins_valid(1) => cond_br252_trueOut_valid,
      ins_ready(0) => cond_br230_falseOut_ready,
      ins_ready(1) => cond_br252_trueOut_ready,
      clk => clk,
      rst => rst,
      outs => mux93_outs,
      outs_valid => mux93_outs_valid,
      outs_ready => mux93_outs_ready
    );

  buffer55 : entity work.oehb(arch) generic map(8)
    port map(
      ins => mux93_outs,
      ins_valid => mux93_outs_valid,
      ins_ready => mux93_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer55_outs,
      outs_valid => buffer55_outs_valid,
      outs_ready => buffer55_outs_ready
    );

  buffer56 : entity work.tehb(arch) generic map(8)
    port map(
      ins => buffer55_outs,
      ins_valid => buffer55_outs_valid,
      ins_ready => buffer55_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer56_outs,
      outs_valid => buffer56_outs_valid,
      outs_ready => buffer56_outs_ready
    );

  fork53 : entity work.handshake_fork(arch) generic map(2, 8)
    port map(
      ins => buffer56_outs,
      ins_valid => buffer56_outs_valid,
      ins_ready => buffer56_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork53_outs_0,
      outs(1) => fork53_outs_1,
      outs_valid(0) => fork53_outs_0_valid,
      outs_valid(1) => fork53_outs_1_valid,
      outs_ready(0) => fork53_outs_0_ready,
      outs_ready(1) => fork53_outs_1_ready
    );

  extsi36 : entity work.extsi(arch) generic map(8, 32)
    port map(
      ins => buffer193_outs,
      ins_valid => buffer193_outs_valid,
      ins_ready => buffer193_outs_ready,
      clk => clk,
      rst => rst,
      outs => extsi36_outs,
      outs_valid => extsi36_outs_valid,
      outs_ready => extsi36_outs_ready
    );

  buffer193 : entity work.tfifo(arch) generic map(1, 8)
    port map(
      ins => fork53_outs_1,
      ins_valid => fork53_outs_1_valid,
      ins_ready => fork53_outs_1_ready,
      clk => clk,
      rst => rst,
      outs => buffer193_outs,
      outs_valid => buffer193_outs_valid,
      outs_ready => buffer193_outs_ready
    );

  mux94 : entity work.mux_dataless(arch) generic map(2, 1)
    port map(
      index => buffer194_outs,
      index_valid => buffer194_outs_valid,
      index_ready => buffer194_outs_ready,
      ins_valid(0) => cond_br226_falseOut_valid,
      ins_valid(1) => cond_br250_trueOut_valid,
      ins_ready(0) => cond_br226_falseOut_ready,
      ins_ready(1) => cond_br250_trueOut_ready,
      clk => clk,
      rst => rst,
      outs_valid => mux94_outs_valid,
      outs_ready => mux94_outs_ready
    );

  buffer194 : entity work.tfifo(arch) generic map(1, 1)
    port map(
      ins => fork52_outs_19,
      ins_valid => fork52_outs_19_valid,
      ins_ready => fork52_outs_19_ready,
      clk => clk,
      rst => rst,
      outs => buffer194_outs,
      outs_valid => buffer194_outs_valid,
      outs_ready => buffer194_outs_ready
    );

  buffer58 : entity work.oehb_dataless(arch)
    port map(
      ins_valid => mux94_outs_valid,
      ins_ready => mux94_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer58_outs_valid,
      outs_ready => buffer58_outs_ready
    );

  buffer59 : entity work.tehb_dataless(arch)
    port map(
      ins_valid => buffer58_outs_valid,
      ins_ready => buffer58_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer59_outs_valid,
      outs_ready => buffer59_outs_ready
    );

  fork54 : entity work.fork_dataless(arch) generic map(2)
    port map(
      ins_valid => buffer59_outs_valid,
      ins_ready => buffer59_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid(0) => fork54_outs_0_valid,
      outs_valid(1) => fork54_outs_1_valid,
      outs_ready(0) => fork54_outs_0_ready,
      outs_ready(1) => fork54_outs_1_ready
    );

  mux95 : entity work.mux(arch) generic map(2, 32, 1)
    port map(
      index => buffer195_outs,
      index_valid => buffer195_outs_valid,
      index_ready => buffer195_outs_ready,
      ins(0) => cond_br225_falseOut,
      ins(1) => cond_br251_trueOut,
      ins_valid(0) => cond_br225_falseOut_valid,
      ins_valid(1) => cond_br251_trueOut_valid,
      ins_ready(0) => cond_br225_falseOut_ready,
      ins_ready(1) => cond_br251_trueOut_ready,
      clk => clk,
      rst => rst,
      outs => mux95_outs,
      outs_valid => mux95_outs_valid,
      outs_ready => mux95_outs_ready
    );

  buffer195 : entity work.tfifo(arch) generic map(1, 1)
    port map(
      ins => fork52_outs_18,
      ins_valid => fork52_outs_18_valid,
      ins_ready => fork52_outs_18_ready,
      clk => clk,
      rst => rst,
      outs => buffer195_outs,
      outs_valid => buffer195_outs_valid,
      outs_ready => buffer195_outs_ready
    );

  buffer60 : entity work.oehb(arch) generic map(32)
    port map(
      ins => mux95_outs,
      ins_valid => mux95_outs_valid,
      ins_ready => mux95_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer60_outs,
      outs_valid => buffer60_outs_valid,
      outs_ready => buffer60_outs_ready
    );

  buffer61 : entity work.tehb(arch) generic map(32)
    port map(
      ins => buffer60_outs,
      ins_valid => buffer60_outs_valid,
      ins_ready => buffer60_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer61_outs,
      outs_valid => buffer61_outs_valid,
      outs_ready => buffer61_outs_ready
    );

  fork55 : entity work.handshake_fork(arch) generic map(2, 32)
    port map(
      ins => buffer61_outs,
      ins_valid => buffer61_outs_valid,
      ins_ready => buffer61_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork55_outs_0,
      outs(1) => fork55_outs_1,
      outs_valid(0) => fork55_outs_0_valid,
      outs_valid(1) => fork55_outs_1_valid,
      outs_ready(0) => fork55_outs_0_ready,
      outs_ready(1) => fork55_outs_1_ready
    );

  mux96 : entity work.mux_dataless(arch) generic map(2, 1)
    port map(
      index => buffer196_outs,
      index_valid => buffer196_outs_valid,
      index_ready => buffer196_outs_ready,
      ins_valid(0) => cond_br223_falseOut_valid,
      ins_valid(1) => cond_br255_trueOut_valid,
      ins_ready(0) => cond_br223_falseOut_ready,
      ins_ready(1) => cond_br255_trueOut_ready,
      clk => clk,
      rst => rst,
      outs_valid => mux96_outs_valid,
      outs_ready => mux96_outs_ready
    );

  buffer196 : entity work.tfifo(arch) generic map(1, 1)
    port map(
      ins => fork52_outs_17,
      ins_valid => fork52_outs_17_valid,
      ins_ready => fork52_outs_17_ready,
      clk => clk,
      rst => rst,
      outs => buffer196_outs,
      outs_valid => buffer196_outs_valid,
      outs_ready => buffer196_outs_ready
    );

  buffer62 : entity work.oehb_dataless(arch)
    port map(
      ins_valid => mux96_outs_valid,
      ins_ready => mux96_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer62_outs_valid,
      outs_ready => buffer62_outs_ready
    );

  buffer63 : entity work.tehb_dataless(arch)
    port map(
      ins_valid => buffer62_outs_valid,
      ins_ready => buffer62_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer63_outs_valid,
      outs_ready => buffer63_outs_ready
    );

  fork56 : entity work.fork_dataless(arch) generic map(2)
    port map(
      ins_valid => buffer63_outs_valid,
      ins_ready => buffer63_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid(0) => fork56_outs_0_valid,
      outs_valid(1) => fork56_outs_1_valid,
      outs_ready(0) => fork56_outs_0_ready,
      outs_ready(1) => fork56_outs_1_ready
    );

  mux97 : entity work.mux(arch) generic map(2, 9, 1)
    port map(
      index => buffer197_outs,
      index_valid => buffer197_outs_valid,
      index_ready => buffer197_outs_ready,
      ins(0) => cond_br220_falseOut,
      ins(1) => cond_br234_trueOut,
      ins_valid(0) => cond_br220_falseOut_valid,
      ins_valid(1) => cond_br234_trueOut_valid,
      ins_ready(0) => cond_br220_falseOut_ready,
      ins_ready(1) => cond_br234_trueOut_ready,
      clk => clk,
      rst => rst,
      outs => mux97_outs,
      outs_valid => mux97_outs_valid,
      outs_ready => mux97_outs_ready
    );

  buffer197 : entity work.tfifo(arch) generic map(1, 1)
    port map(
      ins => fork52_outs_1,
      ins_valid => fork52_outs_1_valid,
      ins_ready => fork52_outs_1_ready,
      clk => clk,
      rst => rst,
      outs => buffer197_outs,
      outs_valid => buffer197_outs_valid,
      outs_ready => buffer197_outs_ready
    );

  buffer64 : entity work.oehb(arch) generic map(9)
    port map(
      ins => mux97_outs,
      ins_valid => mux97_outs_valid,
      ins_ready => mux97_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer64_outs,
      outs_valid => buffer64_outs_valid,
      outs_ready => buffer64_outs_ready
    );

  buffer65 : entity work.tehb(arch) generic map(9)
    port map(
      ins => buffer64_outs,
      ins_valid => buffer64_outs_valid,
      ins_ready => buffer64_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer65_outs,
      outs_valid => buffer65_outs_valid,
      outs_ready => buffer65_outs_ready
    );

  fork57 : entity work.handshake_fork(arch) generic map(2, 9)
    port map(
      ins => buffer65_outs,
      ins_valid => buffer65_outs_valid,
      ins_ready => buffer65_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork57_outs_0,
      outs(1) => fork57_outs_1,
      outs_valid(0) => fork57_outs_0_valid,
      outs_valid(1) => fork57_outs_1_valid,
      outs_ready(0) => fork57_outs_0_ready,
      outs_ready(1) => fork57_outs_1_ready
    );

  extsi37 : entity work.extsi(arch) generic map(9, 32)
    port map(
      ins => buffer198_outs,
      ins_valid => buffer198_outs_valid,
      ins_ready => buffer198_outs_ready,
      clk => clk,
      rst => rst,
      outs => extsi37_outs,
      outs_valid => extsi37_outs_valid,
      outs_ready => extsi37_outs_ready
    );

  buffer198 : entity work.tfifo(arch) generic map(1, 9)
    port map(
      ins => fork57_outs_1,
      ins_valid => fork57_outs_1_valid,
      ins_ready => fork57_outs_1_ready,
      clk => clk,
      rst => rst,
      outs => buffer198_outs,
      outs_valid => buffer198_outs_valid,
      outs_ready => buffer198_outs_ready
    );

  mux98 : entity work.mux(arch) generic map(2, 8, 1)
    port map(
      index => buffer199_outs,
      index_valid => buffer199_outs_valid,
      index_ready => buffer199_outs_ready,
      ins(0) => cond_br212_falseOut,
      ins(1) => cond_br242_trueOut,
      ins_valid(0) => cond_br212_falseOut_valid,
      ins_valid(1) => cond_br242_trueOut_valid,
      ins_ready(0) => cond_br212_falseOut_ready,
      ins_ready(1) => cond_br242_trueOut_ready,
      clk => clk,
      rst => rst,
      outs => mux98_outs,
      outs_valid => mux98_outs_valid,
      outs_ready => mux98_outs_ready
    );

  buffer199 : entity work.tfifo(arch) generic map(1, 1)
    port map(
      ins => fork52_outs_0,
      ins_valid => fork52_outs_0_valid,
      ins_ready => fork52_outs_0_ready,
      clk => clk,
      rst => rst,
      outs => buffer199_outs,
      outs_valid => buffer199_outs_valid,
      outs_ready => buffer199_outs_ready
    );

  buffer67 : entity work.oehb(arch) generic map(8)
    port map(
      ins => mux98_outs,
      ins_valid => mux98_outs_valid,
      ins_ready => mux98_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer67_outs,
      outs_valid => buffer67_outs_valid,
      outs_ready => buffer67_outs_ready
    );

  buffer69 : entity work.tehb(arch) generic map(8)
    port map(
      ins => buffer67_outs,
      ins_valid => buffer67_outs_valid,
      ins_ready => buffer67_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer69_outs,
      outs_valid => buffer69_outs_valid,
      outs_ready => buffer69_outs_ready
    );

  fork58 : entity work.handshake_fork(arch) generic map(2, 8)
    port map(
      ins => buffer69_outs,
      ins_valid => buffer69_outs_valid,
      ins_ready => buffer69_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork58_outs_0,
      outs(1) => fork58_outs_1,
      outs_valid(0) => fork58_outs_0_valid,
      outs_valid(1) => fork58_outs_1_valid,
      outs_ready(0) => fork58_outs_0_ready,
      outs_ready(1) => fork58_outs_1_ready
    );

  extsi38 : entity work.extsi(arch) generic map(8, 32)
    port map(
      ins => buffer200_outs,
      ins_valid => buffer200_outs_valid,
      ins_ready => buffer200_outs_ready,
      clk => clk,
      rst => rst,
      outs => extsi38_outs,
      outs_valid => extsi38_outs_valid,
      outs_ready => extsi38_outs_ready
    );

  buffer200 : entity work.tfifo(arch) generic map(1, 8)
    port map(
      ins => fork58_outs_1,
      ins_valid => fork58_outs_1_valid,
      ins_ready => fork58_outs_1_ready,
      clk => clk,
      rst => rst,
      outs => buffer200_outs,
      outs_valid => buffer200_outs_valid,
      outs_ready => buffer200_outs_ready
    );

  mux99 : entity work.mux(arch) generic map(2, 32, 1)
    port map(
      index => buffer201_outs,
      index_valid => buffer201_outs_valid,
      index_ready => buffer201_outs_ready,
      ins(0) => cond_br211_falseOut,
      ins(1) => cond_br239_trueOut,
      ins_valid(0) => cond_br211_falseOut_valid,
      ins_valid(1) => cond_br239_trueOut_valid,
      ins_ready(0) => cond_br211_falseOut_ready,
      ins_ready(1) => cond_br239_trueOut_ready,
      clk => clk,
      rst => rst,
      outs => mux99_outs,
      outs_valid => mux99_outs_valid,
      outs_ready => mux99_outs_ready
    );

  buffer201 : entity work.tfifo(arch) generic map(1, 1)
    port map(
      ins => fork52_outs_16,
      ins_valid => fork52_outs_16_valid,
      ins_ready => fork52_outs_16_ready,
      clk => clk,
      rst => rst,
      outs => buffer201_outs,
      outs_valid => buffer201_outs_valid,
      outs_ready => buffer201_outs_ready
    );

  buffer70 : entity work.oehb(arch) generic map(32)
    port map(
      ins => mux99_outs,
      ins_valid => mux99_outs_valid,
      ins_ready => mux99_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer70_outs,
      outs_valid => buffer70_outs_valid,
      outs_ready => buffer70_outs_ready
    );

  buffer71 : entity work.tehb(arch) generic map(32)
    port map(
      ins => buffer70_outs,
      ins_valid => buffer70_outs_valid,
      ins_ready => buffer70_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer71_outs,
      outs_valid => buffer71_outs_valid,
      outs_ready => buffer71_outs_ready
    );

  fork59 : entity work.handshake_fork(arch) generic map(2, 32)
    port map(
      ins => buffer71_outs,
      ins_valid => buffer71_outs_valid,
      ins_ready => buffer71_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork59_outs_0,
      outs(1) => fork59_outs_1,
      outs_valid(0) => fork59_outs_0_valid,
      outs_valid(1) => fork59_outs_1_valid,
      outs_ready(0) => fork59_outs_0_ready,
      outs_ready(1) => fork59_outs_1_ready
    );

  mux100 : entity work.mux_dataless(arch) generic map(2, 1)
    port map(
      index => buffer202_outs,
      index_valid => buffer202_outs_valid,
      index_ready => buffer202_outs_ready,
      ins_valid(0) => cond_br206_falseOut_valid,
      ins_valid(1) => cond_br248_trueOut_valid,
      ins_ready(0) => cond_br206_falseOut_ready,
      ins_ready(1) => cond_br248_trueOut_ready,
      clk => clk,
      rst => rst,
      outs_valid => mux100_outs_valid,
      outs_ready => mux100_outs_ready
    );

  buffer202 : entity work.tfifo(arch) generic map(1, 1)
    port map(
      ins => fork52_outs_15,
      ins_valid => fork52_outs_15_valid,
      ins_ready => fork52_outs_15_ready,
      clk => clk,
      rst => rst,
      outs => buffer202_outs,
      outs_valid => buffer202_outs_valid,
      outs_ready => buffer202_outs_ready
    );

  buffer72 : entity work.oehb_dataless(arch)
    port map(
      ins_valid => mux100_outs_valid,
      ins_ready => mux100_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer72_outs_valid,
      outs_ready => buffer72_outs_ready
    );

  buffer73 : entity work.tehb_dataless(arch)
    port map(
      ins_valid => buffer72_outs_valid,
      ins_ready => buffer72_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer73_outs_valid,
      outs_ready => buffer73_outs_ready
    );

  fork60 : entity work.fork_dataless(arch) generic map(2)
    port map(
      ins_valid => buffer73_outs_valid,
      ins_ready => buffer73_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid(0) => fork60_outs_0_valid,
      outs_valid(1) => fork60_outs_1_valid,
      outs_ready(0) => fork60_outs_0_ready,
      outs_ready(1) => fork60_outs_1_ready
    );

  mux101 : entity work.mux_dataless(arch) generic map(2, 1)
    port map(
      index => buffer203_outs,
      index_valid => buffer203_outs_valid,
      index_ready => buffer203_outs_ready,
      ins_valid(0) => cond_br219_falseOut_valid,
      ins_valid(1) => cond_br237_trueOut_valid,
      ins_ready(0) => cond_br219_falseOut_ready,
      ins_ready(1) => cond_br237_trueOut_ready,
      clk => clk,
      rst => rst,
      outs_valid => mux101_outs_valid,
      outs_ready => mux101_outs_ready
    );

  buffer203 : entity work.tfifo(arch) generic map(1, 1)
    port map(
      ins => fork52_outs_14,
      ins_valid => fork52_outs_14_valid,
      ins_ready => fork52_outs_14_ready,
      clk => clk,
      rst => rst,
      outs => buffer203_outs,
      outs_valid => buffer203_outs_valid,
      outs_ready => buffer203_outs_ready
    );

  buffer74 : entity work.oehb_dataless(arch)
    port map(
      ins_valid => mux101_outs_valid,
      ins_ready => mux101_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer74_outs_valid,
      outs_ready => buffer74_outs_ready
    );

  buffer75 : entity work.tehb_dataless(arch)
    port map(
      ins_valid => buffer74_outs_valid,
      ins_ready => buffer74_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer75_outs_valid,
      outs_ready => buffer75_outs_ready
    );

  fork61 : entity work.fork_dataless(arch) generic map(2)
    port map(
      ins_valid => buffer75_outs_valid,
      ins_ready => buffer75_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid(0) => fork61_outs_0_valid,
      outs_valid(1) => fork61_outs_1_valid,
      outs_ready(0) => fork61_outs_0_ready,
      outs_ready(1) => fork61_outs_1_ready
    );

  mux102 : entity work.mux_dataless(arch) generic map(2, 1)
    port map(
      index => buffer204_outs,
      index_valid => buffer204_outs_valid,
      index_ready => buffer204_outs_ready,
      ins_valid(0) => cond_br214_falseOut_valid,
      ins_valid(1) => cond_br236_trueOut_valid,
      ins_ready(0) => cond_br214_falseOut_ready,
      ins_ready(1) => cond_br236_trueOut_ready,
      clk => clk,
      rst => rst,
      outs_valid => mux102_outs_valid,
      outs_ready => mux102_outs_ready
    );

  buffer204 : entity work.tfifo(arch) generic map(1, 1)
    port map(
      ins => fork52_outs_13,
      ins_valid => fork52_outs_13_valid,
      ins_ready => fork52_outs_13_ready,
      clk => clk,
      rst => rst,
      outs => buffer204_outs,
      outs_valid => buffer204_outs_valid,
      outs_ready => buffer204_outs_ready
    );

  buffer76 : entity work.oehb_dataless(arch)
    port map(
      ins_valid => mux102_outs_valid,
      ins_ready => mux102_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer76_outs_valid,
      outs_ready => buffer76_outs_ready
    );

  buffer77 : entity work.tehb_dataless(arch)
    port map(
      ins_valid => buffer76_outs_valid,
      ins_ready => buffer76_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer77_outs_valid,
      outs_ready => buffer77_outs_ready
    );

  fork62 : entity work.fork_dataless(arch) generic map(2)
    port map(
      ins_valid => buffer77_outs_valid,
      ins_ready => buffer77_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid(0) => fork62_outs_0_valid,
      outs_valid(1) => fork62_outs_1_valid,
      outs_ready(0) => fork62_outs_0_ready,
      outs_ready(1) => fork62_outs_1_ready
    );

  mux103 : entity work.mux(arch) generic map(2, 32, 1)
    port map(
      index => buffer205_outs,
      index_valid => buffer205_outs_valid,
      index_ready => buffer205_outs_ready,
      ins(0) => cond_br227_falseOut,
      ins(1) => cond_br256_trueOut,
      ins_valid(0) => cond_br227_falseOut_valid,
      ins_valid(1) => cond_br256_trueOut_valid,
      ins_ready(0) => cond_br227_falseOut_ready,
      ins_ready(1) => cond_br256_trueOut_ready,
      clk => clk,
      rst => rst,
      outs => mux103_outs,
      outs_valid => mux103_outs_valid,
      outs_ready => mux103_outs_ready
    );

  buffer205 : entity work.tfifo(arch) generic map(1, 1)
    port map(
      ins => fork52_outs_12,
      ins_valid => fork52_outs_12_valid,
      ins_ready => fork52_outs_12_ready,
      clk => clk,
      rst => rst,
      outs => buffer205_outs,
      outs_valid => buffer205_outs_valid,
      outs_ready => buffer205_outs_ready
    );

  buffer78 : entity work.oehb(arch) generic map(32)
    port map(
      ins => mux103_outs,
      ins_valid => mux103_outs_valid,
      ins_ready => mux103_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer78_outs,
      outs_valid => buffer78_outs_valid,
      outs_ready => buffer78_outs_ready
    );

  buffer79 : entity work.tehb(arch) generic map(32)
    port map(
      ins => buffer78_outs,
      ins_valid => buffer78_outs_valid,
      ins_ready => buffer78_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer79_outs,
      outs_valid => buffer79_outs_valid,
      outs_ready => buffer79_outs_ready
    );

  fork63 : entity work.handshake_fork(arch) generic map(2, 32)
    port map(
      ins => buffer79_outs,
      ins_valid => buffer79_outs_valid,
      ins_ready => buffer79_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork63_outs_0,
      outs(1) => fork63_outs_1,
      outs_valid(0) => fork63_outs_0_valid,
      outs_valid(1) => fork63_outs_1_valid,
      outs_ready(0) => fork63_outs_0_ready,
      outs_ready(1) => fork63_outs_1_ready
    );

  mux104 : entity work.mux_dataless(arch) generic map(2, 1)
    port map(
      index => buffer206_outs,
      index_valid => buffer206_outs_valid,
      index_ready => buffer206_outs_ready,
      ins_valid(0) => cond_br229_falseOut_valid,
      ins_valid(1) => cond_br238_trueOut_valid,
      ins_ready(0) => cond_br229_falseOut_ready,
      ins_ready(1) => cond_br238_trueOut_ready,
      clk => clk,
      rst => rst,
      outs_valid => mux104_outs_valid,
      outs_ready => mux104_outs_ready
    );

  buffer206 : entity work.tfifo(arch) generic map(1, 1)
    port map(
      ins => fork52_outs_11,
      ins_valid => fork52_outs_11_valid,
      ins_ready => fork52_outs_11_ready,
      clk => clk,
      rst => rst,
      outs => buffer206_outs,
      outs_valid => buffer206_outs_valid,
      outs_ready => buffer206_outs_ready
    );

  buffer80 : entity work.oehb_dataless(arch)
    port map(
      ins_valid => mux104_outs_valid,
      ins_ready => mux104_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer80_outs_valid,
      outs_ready => buffer80_outs_ready
    );

  buffer81 : entity work.tehb_dataless(arch)
    port map(
      ins_valid => buffer80_outs_valid,
      ins_ready => buffer80_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer81_outs_valid,
      outs_ready => buffer81_outs_ready
    );

  fork64 : entity work.fork_dataless(arch) generic map(2)
    port map(
      ins_valid => buffer81_outs_valid,
      ins_ready => buffer81_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid(0) => fork64_outs_0_valid,
      outs_valid(1) => fork64_outs_1_valid,
      outs_ready(0) => fork64_outs_0_ready,
      outs_ready(1) => fork64_outs_1_ready
    );

  mux105 : entity work.mux_dataless(arch) generic map(2, 1)
    port map(
      index => buffer207_outs,
      index_valid => buffer207_outs_valid,
      index_ready => buffer207_outs_ready,
      ins_valid(0) => cond_br208_falseOut_valid,
      ins_valid(1) => cond_br240_trueOut_valid,
      ins_ready(0) => cond_br208_falseOut_ready,
      ins_ready(1) => cond_br240_trueOut_ready,
      clk => clk,
      rst => rst,
      outs_valid => mux105_outs_valid,
      outs_ready => mux105_outs_ready
    );

  buffer207 : entity work.tfifo(arch) generic map(1, 1)
    port map(
      ins => fork52_outs_10,
      ins_valid => fork52_outs_10_valid,
      ins_ready => fork52_outs_10_ready,
      clk => clk,
      rst => rst,
      outs => buffer207_outs,
      outs_valid => buffer207_outs_valid,
      outs_ready => buffer207_outs_ready
    );

  buffer82 : entity work.oehb_dataless(arch)
    port map(
      ins_valid => mux105_outs_valid,
      ins_ready => mux105_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer82_outs_valid,
      outs_ready => buffer82_outs_ready
    );

  buffer83 : entity work.tehb_dataless(arch)
    port map(
      ins_valid => buffer82_outs_valid,
      ins_ready => buffer82_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer83_outs_valid,
      outs_ready => buffer83_outs_ready
    );

  fork65 : entity work.fork_dataless(arch) generic map(2)
    port map(
      ins_valid => buffer83_outs_valid,
      ins_ready => buffer83_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid(0) => fork65_outs_0_valid,
      outs_valid(1) => fork65_outs_1_valid,
      outs_ready(0) => fork65_outs_0_ready,
      outs_ready(1) => fork65_outs_1_ready
    );

  mux106 : entity work.mux_dataless(arch) generic map(2, 1)
    port map(
      index => fork52_outs_9,
      index_valid => fork52_outs_9_valid,
      index_ready => fork52_outs_9_ready,
      ins_valid(0) => cond_br210_falseOut_valid,
      ins_valid(1) => cond_br241_trueOut_valid,
      ins_ready(0) => cond_br210_falseOut_ready,
      ins_ready(1) => cond_br241_trueOut_ready,
      clk => clk,
      rst => rst,
      outs_valid => mux106_outs_valid,
      outs_ready => mux106_outs_ready
    );

  buffer84 : entity work.oehb_dataless(arch)
    port map(
      ins_valid => mux106_outs_valid,
      ins_ready => mux106_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer84_outs_valid,
      outs_ready => buffer84_outs_ready
    );

  buffer85 : entity work.tehb_dataless(arch)
    port map(
      ins_valid => buffer84_outs_valid,
      ins_ready => buffer84_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer85_outs_valid,
      outs_ready => buffer85_outs_ready
    );

  fork66 : entity work.fork_dataless(arch) generic map(2)
    port map(
      ins_valid => buffer85_outs_valid,
      ins_ready => buffer85_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid(0) => fork66_outs_0_valid,
      outs_valid(1) => fork66_outs_1_valid,
      outs_ready(0) => fork66_outs_0_ready,
      outs_ready(1) => fork66_outs_1_ready
    );

  mux107 : entity work.mux_dataless(arch) generic map(2, 1)
    port map(
      index => buffer209_outs,
      index_valid => buffer209_outs_valid,
      index_ready => buffer209_outs_ready,
      ins_valid(0) => cond_br221_falseOut_valid,
      ins_valid(1) => cond_br247_trueOut_valid,
      ins_ready(0) => cond_br221_falseOut_ready,
      ins_ready(1) => cond_br247_trueOut_ready,
      clk => clk,
      rst => rst,
      outs_valid => mux107_outs_valid,
      outs_ready => mux107_outs_ready
    );

  buffer209 : entity work.tfifo(arch) generic map(1, 1)
    port map(
      ins => fork52_outs_8,
      ins_valid => fork52_outs_8_valid,
      ins_ready => fork52_outs_8_ready,
      clk => clk,
      rst => rst,
      outs => buffer209_outs,
      outs_valid => buffer209_outs_valid,
      outs_ready => buffer209_outs_ready
    );

  buffer86 : entity work.oehb_dataless(arch)
    port map(
      ins_valid => mux107_outs_valid,
      ins_ready => mux107_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer86_outs_valid,
      outs_ready => buffer86_outs_ready
    );

  buffer87 : entity work.tehb_dataless(arch)
    port map(
      ins_valid => buffer86_outs_valid,
      ins_ready => buffer86_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer87_outs_valid,
      outs_ready => buffer87_outs_ready
    );

  fork67 : entity work.fork_dataless(arch) generic map(2)
    port map(
      ins_valid => buffer87_outs_valid,
      ins_ready => buffer87_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid(0) => fork67_outs_0_valid,
      outs_valid(1) => fork67_outs_1_valid,
      outs_ready(0) => fork67_outs_0_ready,
      outs_ready(1) => fork67_outs_1_ready
    );

  mux108 : entity work.mux_dataless(arch) generic map(2, 1)
    port map(
      index => buffer210_outs,
      index_valid => buffer210_outs_valid,
      index_ready => buffer210_outs_ready,
      ins_valid(0) => cond_br231_falseOut_valid,
      ins_valid(1) => cond_br253_trueOut_valid,
      ins_ready(0) => cond_br231_falseOut_ready,
      ins_ready(1) => cond_br253_trueOut_ready,
      clk => clk,
      rst => rst,
      outs_valid => mux108_outs_valid,
      outs_ready => mux108_outs_ready
    );

  buffer210 : entity work.tfifo(arch) generic map(1, 1)
    port map(
      ins => fork52_outs_7,
      ins_valid => fork52_outs_7_valid,
      ins_ready => fork52_outs_7_ready,
      clk => clk,
      rst => rst,
      outs => buffer210_outs,
      outs_valid => buffer210_outs_valid,
      outs_ready => buffer210_outs_ready
    );

  buffer88 : entity work.oehb_dataless(arch)
    port map(
      ins_valid => mux108_outs_valid,
      ins_ready => mux108_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer88_outs_valid,
      outs_ready => buffer88_outs_ready
    );

  buffer89 : entity work.tehb_dataless(arch)
    port map(
      ins_valid => buffer88_outs_valid,
      ins_ready => buffer88_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer89_outs_valid,
      outs_ready => buffer89_outs_ready
    );

  fork68 : entity work.fork_dataless(arch) generic map(2)
    port map(
      ins_valid => buffer89_outs_valid,
      ins_ready => buffer89_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid(0) => fork68_outs_0_valid,
      outs_valid(1) => fork68_outs_1_valid,
      outs_ready(0) => fork68_outs_0_ready,
      outs_ready(1) => fork68_outs_1_ready
    );

  mux109 : entity work.mux(arch) generic map(2, 32, 1)
    port map(
      index => buffer211_outs,
      index_valid => buffer211_outs_valid,
      index_ready => buffer211_outs_ready,
      ins(0) => cond_br232_falseOut,
      ins(1) => cond_br254_trueOut,
      ins_valid(0) => cond_br232_falseOut_valid,
      ins_valid(1) => cond_br254_trueOut_valid,
      ins_ready(0) => cond_br232_falseOut_ready,
      ins_ready(1) => cond_br254_trueOut_ready,
      clk => clk,
      rst => rst,
      outs => mux109_outs,
      outs_valid => mux109_outs_valid,
      outs_ready => mux109_outs_ready
    );

  buffer211 : entity work.tfifo(arch) generic map(1, 1)
    port map(
      ins => fork52_outs_6,
      ins_valid => fork52_outs_6_valid,
      ins_ready => fork52_outs_6_ready,
      clk => clk,
      rst => rst,
      outs => buffer211_outs,
      outs_valid => buffer211_outs_valid,
      outs_ready => buffer211_outs_ready
    );

  buffer90 : entity work.oehb(arch) generic map(32)
    port map(
      ins => mux109_outs,
      ins_valid => mux109_outs_valid,
      ins_ready => mux109_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer90_outs,
      outs_valid => buffer90_outs_valid,
      outs_ready => buffer90_outs_ready
    );

  buffer91 : entity work.tehb(arch) generic map(32)
    port map(
      ins => buffer90_outs,
      ins_valid => buffer90_outs_valid,
      ins_ready => buffer90_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer91_outs,
      outs_valid => buffer91_outs_valid,
      outs_ready => buffer91_outs_ready
    );

  fork69 : entity work.handshake_fork(arch) generic map(2, 32)
    port map(
      ins => buffer91_outs,
      ins_valid => buffer91_outs_valid,
      ins_ready => buffer91_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork69_outs_0,
      outs(1) => fork69_outs_1,
      outs_valid(0) => fork69_outs_0_valid,
      outs_valid(1) => fork69_outs_1_valid,
      outs_ready(0) => fork69_outs_0_ready,
      outs_ready(1) => fork69_outs_1_ready
    );

  mux110 : entity work.mux(arch) generic map(2, 32, 1)
    port map(
      index => buffer212_outs,
      index_valid => buffer212_outs_valid,
      index_ready => buffer212_outs_ready,
      ins(0) => cond_br224_falseOut,
      ins(1) => cond_br235_trueOut,
      ins_valid(0) => cond_br224_falseOut_valid,
      ins_valid(1) => cond_br235_trueOut_valid,
      ins_ready(0) => cond_br224_falseOut_ready,
      ins_ready(1) => cond_br235_trueOut_ready,
      clk => clk,
      rst => rst,
      outs => mux110_outs,
      outs_valid => mux110_outs_valid,
      outs_ready => mux110_outs_ready
    );

  buffer212 : entity work.tfifo(arch) generic map(1, 1)
    port map(
      ins => fork52_outs_5,
      ins_valid => fork52_outs_5_valid,
      ins_ready => fork52_outs_5_ready,
      clk => clk,
      rst => rst,
      outs => buffer212_outs,
      outs_valid => buffer212_outs_valid,
      outs_ready => buffer212_outs_ready
    );

  buffer92 : entity work.oehb(arch) generic map(32)
    port map(
      ins => mux110_outs,
      ins_valid => mux110_outs_valid,
      ins_ready => mux110_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer92_outs,
      outs_valid => buffer92_outs_valid,
      outs_ready => buffer92_outs_ready
    );

  buffer93 : entity work.tehb(arch) generic map(32)
    port map(
      ins => buffer92_outs,
      ins_valid => buffer92_outs_valid,
      ins_ready => buffer92_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer93_outs,
      outs_valid => buffer93_outs_valid,
      outs_ready => buffer93_outs_ready
    );

  fork70 : entity work.handshake_fork(arch) generic map(2, 32)
    port map(
      ins => buffer93_outs,
      ins_valid => buffer93_outs_valid,
      ins_ready => buffer93_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork70_outs_0,
      outs(1) => fork70_outs_1,
      outs_valid(0) => fork70_outs_0_valid,
      outs_valid(1) => fork70_outs_1_valid,
      outs_ready(0) => fork70_outs_0_ready,
      outs_ready(1) => fork70_outs_1_ready
    );

  mux111 : entity work.mux_dataless(arch) generic map(2, 1)
    port map(
      index => buffer213_outs,
      index_valid => buffer213_outs_valid,
      index_ready => buffer213_outs_ready,
      ins_valid(0) => cond_br216_falseOut_valid,
      ins_valid(1) => cond_br243_trueOut_valid,
      ins_ready(0) => cond_br216_falseOut_ready,
      ins_ready(1) => cond_br243_trueOut_ready,
      clk => clk,
      rst => rst,
      outs_valid => mux111_outs_valid,
      outs_ready => mux111_outs_ready
    );

  buffer213 : entity work.tfifo(arch) generic map(1, 1)
    port map(
      ins => fork52_outs_4,
      ins_valid => fork52_outs_4_valid,
      ins_ready => fork52_outs_4_ready,
      clk => clk,
      rst => rst,
      outs => buffer213_outs,
      outs_valid => buffer213_outs_valid,
      outs_ready => buffer213_outs_ready
    );

  buffer94 : entity work.oehb_dataless(arch)
    port map(
      ins_valid => mux111_outs_valid,
      ins_ready => mux111_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer94_outs_valid,
      outs_ready => buffer94_outs_ready
    );

  buffer95 : entity work.tehb_dataless(arch)
    port map(
      ins_valid => buffer94_outs_valid,
      ins_ready => buffer94_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer95_outs_valid,
      outs_ready => buffer95_outs_ready
    );

  fork71 : entity work.fork_dataless(arch) generic map(2)
    port map(
      ins_valid => buffer95_outs_valid,
      ins_ready => buffer95_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid(0) => fork71_outs_0_valid,
      outs_valid(1) => fork71_outs_1_valid,
      outs_ready(0) => fork71_outs_0_ready,
      outs_ready(1) => fork71_outs_1_ready
    );

  mux112 : entity work.mux_dataless(arch) generic map(2, 1)
    port map(
      index => buffer214_outs,
      index_valid => buffer214_outs_valid,
      index_ready => buffer214_outs_ready,
      ins_valid(0) => cond_br215_falseOut_valid,
      ins_valid(1) => cond_br245_trueOut_valid,
      ins_ready(0) => cond_br215_falseOut_ready,
      ins_ready(1) => cond_br245_trueOut_ready,
      clk => clk,
      rst => rst,
      outs_valid => mux112_outs_valid,
      outs_ready => mux112_outs_ready
    );

  buffer214 : entity work.tfifo(arch) generic map(1, 1)
    port map(
      ins => fork52_outs_3,
      ins_valid => fork52_outs_3_valid,
      ins_ready => fork52_outs_3_ready,
      clk => clk,
      rst => rst,
      outs => buffer214_outs,
      outs_valid => buffer214_outs_valid,
      outs_ready => buffer214_outs_ready
    );

  buffer96 : entity work.oehb_dataless(arch)
    port map(
      ins_valid => mux112_outs_valid,
      ins_ready => mux112_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer96_outs_valid,
      outs_ready => buffer96_outs_ready
    );

  buffer97 : entity work.tehb_dataless(arch)
    port map(
      ins_valid => buffer96_outs_valid,
      ins_ready => buffer96_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer97_outs_valid,
      outs_ready => buffer97_outs_ready
    );

  fork72 : entity work.fork_dataless(arch) generic map(2)
    port map(
      ins_valid => buffer97_outs_valid,
      ins_ready => buffer97_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid(0) => fork72_outs_0_valid,
      outs_valid(1) => fork72_outs_1_valid,
      outs_ready(0) => fork72_outs_0_ready,
      outs_ready(1) => fork72_outs_1_ready
    );

  unbundle7 : entity work.unbundle(arch) generic map(32)
    port map(
      ins => fork81_outs_1,
      ins_valid => fork81_outs_1_valid,
      ins_ready => fork81_outs_1_ready,
      clk => clk,
      rst => rst,
      outs_valid => unbundle7_outs_0_valid,
      outs_ready => unbundle7_outs_0_ready,
      outs => unbundle7_outs_1
    );

  mux3 : entity work.mux(arch) generic map(2, 8, 1)
    port map(
      index => fork75_outs_1,
      index_valid => fork75_outs_1_valid,
      index_ready => fork75_outs_1_ready,
      ins(0) => extsi19_outs,
      ins(1) => cond_br7_trueOut,
      ins_valid(0) => extsi19_outs_valid,
      ins_valid(1) => cond_br7_trueOut_valid,
      ins_ready(0) => extsi19_outs_ready,
      ins_ready(1) => cond_br7_trueOut_ready,
      clk => clk,
      rst => rst,
      outs => mux3_outs,
      outs_valid => mux3_outs_valid,
      outs_ready => mux3_outs_ready
    );

  buffer98 : entity work.oehb(arch) generic map(8)
    port map(
      ins => mux3_outs,
      ins_valid => mux3_outs_valid,
      ins_ready => mux3_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer98_outs,
      outs_valid => buffer98_outs_valid,
      outs_ready => buffer98_outs_ready
    );

  buffer99 : entity work.tehb(arch) generic map(8)
    port map(
      ins => buffer98_outs,
      ins_valid => buffer98_outs_valid,
      ins_ready => buffer98_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer99_outs,
      outs_valid => buffer99_outs_valid,
      outs_ready => buffer99_outs_ready
    );

  fork73 : entity work.handshake_fork(arch) generic map(4, 8)
    port map(
      ins => buffer99_outs,
      ins_valid => buffer99_outs_valid,
      ins_ready => buffer99_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork73_outs_0,
      outs(1) => fork73_outs_1,
      outs(2) => fork73_outs_2,
      outs(3) => fork73_outs_3,
      outs_valid(0) => fork73_outs_0_valid,
      outs_valid(1) => fork73_outs_1_valid,
      outs_valid(2) => fork73_outs_2_valid,
      outs_valid(3) => fork73_outs_3_valid,
      outs_ready(0) => fork73_outs_0_ready,
      outs_ready(1) => fork73_outs_1_ready,
      outs_ready(2) => fork73_outs_2_ready,
      outs_ready(3) => fork73_outs_3_ready
    );

  extsi39 : entity work.extsi(arch) generic map(8, 9)
    port map(
      ins => fork73_outs_0,
      ins_valid => fork73_outs_0_valid,
      ins_ready => fork73_outs_0_ready,
      clk => clk,
      rst => rst,
      outs => extsi39_outs,
      outs_valid => extsi39_outs_valid,
      outs_ready => extsi39_outs_ready
    );

  extsi40 : entity work.extsi(arch) generic map(8, 32)
    port map(
      ins => buffer218_outs,
      ins_valid => buffer218_outs_valid,
      ins_ready => buffer218_outs_ready,
      clk => clk,
      rst => rst,
      outs => extsi40_outs,
      outs_valid => extsi40_outs_valid,
      outs_ready => extsi40_outs_ready
    );

  buffer218 : entity work.tfifo(arch) generic map(1, 8)
    port map(
      ins => fork73_outs_3,
      ins_valid => fork73_outs_3_valid,
      ins_ready => fork73_outs_3_ready,
      clk => clk,
      rst => rst,
      outs => buffer218_outs,
      outs_valid => buffer218_outs_valid,
      outs_ready => buffer218_outs_ready
    );

  fork74 : entity work.handshake_fork(arch) generic map(6, 32)
    port map(
      ins => extsi40_outs,
      ins_valid => extsi40_outs_valid,
      ins_ready => extsi40_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork74_outs_0,
      outs(1) => fork74_outs_1,
      outs(2) => fork74_outs_2,
      outs(3) => fork74_outs_3,
      outs(4) => fork74_outs_4,
      outs(5) => fork74_outs_5,
      outs_valid(0) => fork74_outs_0_valid,
      outs_valid(1) => fork74_outs_1_valid,
      outs_valid(2) => fork74_outs_2_valid,
      outs_valid(3) => fork74_outs_3_valid,
      outs_valid(4) => fork74_outs_4_valid,
      outs_valid(5) => fork74_outs_5_valid,
      outs_ready(0) => fork74_outs_0_ready,
      outs_ready(1) => fork74_outs_1_ready,
      outs_ready(2) => fork74_outs_2_ready,
      outs_ready(3) => fork74_outs_3_ready,
      outs_ready(4) => fork74_outs_4_ready,
      outs_ready(5) => fork74_outs_5_ready
    );

  mux4 : entity work.mux(arch) generic map(2, 3, 1)
    port map(
      index => fork75_outs_0,
      index_valid => fork75_outs_0_valid,
      index_ready => fork75_outs_0_ready,
      ins(0) => cond_br4_falseOut,
      ins(1) => cond_br8_trueOut,
      ins_valid(0) => cond_br4_falseOut_valid,
      ins_valid(1) => cond_br8_trueOut_valid,
      ins_ready(0) => cond_br4_falseOut_ready,
      ins_ready(1) => cond_br8_trueOut_ready,
      clk => clk,
      rst => rst,
      outs => mux4_outs,
      outs_valid => mux4_outs_valid,
      outs_ready => mux4_outs_ready
    );

  control_merge2 : entity work.control_merge_dataless(arch) generic map(2, 1)
    port map(
      ins_valid(0) => cond_br5_falseOut_valid,
      ins_valid(1) => cond_br9_trueOut_valid,
      ins_ready(0) => cond_br5_falseOut_ready,
      ins_ready(1) => cond_br9_trueOut_ready,
      clk => clk,
      rst => rst,
      outs_valid => control_merge2_outs_valid,
      outs_ready => control_merge2_outs_ready,
      index => control_merge2_index,
      index_valid => control_merge2_index_valid,
      index_ready => control_merge2_index_ready
    );

  fork75 : entity work.handshake_fork(arch) generic map(2, 1)
    port map(
      ins => control_merge2_index,
      ins_valid => control_merge2_index_valid,
      ins_ready => control_merge2_index_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork75_outs_0,
      outs(1) => fork75_outs_1,
      outs_valid(0) => fork75_outs_0_valid,
      outs_valid(1) => fork75_outs_1_valid,
      outs_ready(0) => fork75_outs_0_ready,
      outs_ready(1) => fork75_outs_1_ready
    );

  fork76 : entity work.fork_dataless(arch) generic map(2)
    port map(
      ins_valid => control_merge2_outs_valid,
      ins_ready => control_merge2_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid(0) => fork76_outs_0_valid,
      outs_valid(1) => fork76_outs_1_valid,
      outs_ready(0) => fork76_outs_0_ready,
      outs_ready(1) => fork76_outs_1_ready
    );

  constant20 : entity work.handshake_constant_2(arch) generic map(2)
    port map(
      ctrl_valid => fork76_outs_0_valid,
      ctrl_ready => fork76_outs_0_ready,
      clk => clk,
      rst => rst,
      outs => constant20_outs,
      outs_valid => constant20_outs_valid,
      outs_ready => constant20_outs_ready
    );

  extsi14 : entity work.extsi(arch) generic map(2, 32)
    port map(
      ins => constant20_outs,
      ins_valid => constant20_outs_valid,
      ins_ready => constant20_outs_ready,
      clk => clk,
      rst => rst,
      outs => extsi14_outs,
      outs_valid => extsi14_outs_valid,
      outs_ready => extsi14_outs_ready
    );

  source3 : entity work.source(arch)
    port map(
      clk => clk,
      rst => rst,
      outs_valid => source3_outs_valid,
      outs_ready => source3_outs_ready
    );

  constant25 : entity work.handshake_constant_4(arch) generic map(8)
    port map(
      ctrl_valid => source3_outs_valid,
      ctrl_ready => source3_outs_ready,
      clk => clk,
      rst => rst,
      outs => constant25_outs,
      outs_valid => constant25_outs_valid,
      outs_ready => constant25_outs_ready
    );

  extsi41 : entity work.extsi(arch) generic map(8, 9)
    port map(
      ins => constant25_outs,
      ins_valid => constant25_outs_valid,
      ins_ready => constant25_outs_ready,
      clk => clk,
      rst => rst,
      outs => extsi41_outs,
      outs_valid => extsi41_outs_valid,
      outs_ready => extsi41_outs_ready
    );

  source4 : entity work.source(arch)
    port map(
      clk => clk,
      rst => rst,
      outs_valid => source4_outs_valid,
      outs_ready => source4_outs_ready
    );

  constant28 : entity work.handshake_constant_2(arch) generic map(2)
    port map(
      ctrl_valid => source4_outs_valid,
      ctrl_ready => source4_outs_ready,
      clk => clk,
      rst => rst,
      outs => constant28_outs,
      outs_valid => constant28_outs_valid,
      outs_ready => constant28_outs_ready
    );

  extsi42 : entity work.extsi(arch) generic map(2, 9)
    port map(
      ins => constant28_outs,
      ins_valid => constant28_outs_valid,
      ins_ready => constant28_outs_ready,
      clk => clk,
      rst => rst,
      outs => extsi42_outs,
      outs_valid => extsi42_outs_valid,
      outs_ready => extsi42_outs_ready
    );

  gate8 : entity work.gate(arch) generic map(2, 32)
    port map(
      ins(0) => buffer220_outs,
      ins_valid(0) => buffer220_outs_valid,
      ins_valid(1) => fork62_outs_0_valid,
      ins_ready(0) => buffer220_outs_ready,
      ins_ready(1) => fork62_outs_0_ready,
      clk => clk,
      rst => rst,
      outs => gate8_outs,
      outs_valid => gate8_outs_valid,
      outs_ready => gate8_outs_ready
    );

  buffer220 : entity work.tfifo(arch) generic map(1, 32)
    port map(
      ins => fork74_outs_0,
      ins_valid => fork74_outs_0_valid,
      ins_ready => fork74_outs_0_ready,
      clk => clk,
      rst => rst,
      outs => buffer220_outs,
      outs_valid => buffer220_outs_valid,
      outs_ready => buffer220_outs_ready
    );

  fork77 : entity work.handshake_fork(arch) generic map(2, 32)
    port map(
      ins => gate8_outs,
      ins_valid => gate8_outs_valid,
      ins_ready => gate8_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork77_outs_0,
      outs(1) => fork77_outs_1,
      outs_valid(0) => fork77_outs_0_valid,
      outs_valid(1) => fork77_outs_1_valid,
      outs_ready(0) => fork77_outs_0_ready,
      outs_ready(1) => fork77_outs_1_ready
    );

  cmpi11 : entity work.handshake_cmpi_0(arch) generic map(32)
    port map(
      lhs => fork77_outs_1,
      lhs_valid => fork77_outs_1_valid,
      lhs_ready => fork77_outs_1_ready,
      rhs => extsi38_outs,
      rhs_valid => extsi38_outs_valid,
      rhs_ready => extsi38_outs_ready,
      clk => clk,
      rst => rst,
      result => cmpi11_result,
      result_valid => cmpi11_result_valid,
      result_ready => cmpi11_result_ready
    );

  fork78 : entity work.handshake_fork(arch) generic map(2, 1)
    port map(
      ins => cmpi11_result,
      ins_valid => cmpi11_result_valid,
      ins_ready => cmpi11_result_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork78_outs_0,
      outs(1) => fork78_outs_1,
      outs_valid(0) => fork78_outs_0_valid,
      outs_valid(1) => fork78_outs_1_valid,
      outs_ready(0) => fork78_outs_0_ready,
      outs_ready(1) => fork78_outs_1_ready
    );

  cmpi12 : entity work.handshake_cmpi_0(arch) generic map(32)
    port map(
      lhs => fork77_outs_0,
      lhs_valid => fork77_outs_0_valid,
      lhs_ready => fork77_outs_0_ready,
      rhs => buffer223_outs,
      rhs_valid => buffer223_outs_valid,
      rhs_ready => buffer223_outs_ready,
      clk => clk,
      rst => rst,
      result => cmpi12_result,
      result_valid => cmpi12_result_valid,
      result_ready => cmpi12_result_ready
    );

  buffer223 : entity work.tfifo(arch) generic map(1, 32)
    port map(
      ins => fork59_outs_0,
      ins_valid => fork59_outs_0_valid,
      ins_ready => fork59_outs_0_ready,
      clk => clk,
      rst => rst,
      outs => buffer223_outs,
      outs_valid => buffer223_outs_valid,
      outs_ready => buffer223_outs_ready
    );

  fork79 : entity work.handshake_fork(arch) generic map(2, 1)
    port map(
      ins => cmpi12_result,
      ins_valid => cmpi12_result_valid,
      ins_ready => cmpi12_result_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork79_outs_0,
      outs(1) => fork79_outs_1,
      outs_valid(0) => fork79_outs_0_valid,
      outs_valid(1) => fork79_outs_1_valid,
      outs_ready(0) => fork79_outs_0_ready,
      outs_ready(1) => fork79_outs_1_ready
    );

  buffer8 : entity work.tfifo(arch) generic map(1, 8)
    port map(
      ins => fork73_outs_2,
      ins_valid => fork73_outs_2_valid,
      ins_ready => fork73_outs_2_ready,
      clk => clk,
      rst => rst,
      outs => buffer8_outs,
      outs_valid => buffer8_outs_valid,
      outs_ready => buffer8_outs_ready
    );

  fork80 : entity work.handshake_fork(arch) generic map(2, 8)
    port map(
      ins => buffer8_outs,
      ins_valid => buffer8_outs_valid,
      ins_ready => buffer8_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork80_outs_0,
      outs(1) => fork80_outs_1,
      outs_valid(0) => fork80_outs_0_valid,
      outs_valid(1) => fork80_outs_1_valid,
      outs_ready(0) => fork80_outs_0_ready,
      outs_ready(1) => fork80_outs_1_ready
    );

  extsi43 : entity work.extsi(arch) generic map(8, 32)
    port map(
      ins => buffer225_outs,
      ins_valid => buffer225_outs_valid,
      ins_ready => buffer225_outs_ready,
      clk => clk,
      rst => rst,
      outs => extsi43_outs,
      outs_valid => extsi43_outs_valid,
      outs_ready => extsi43_outs_ready
    );

  buffer225 : entity work.tfifo(arch) generic map(1, 8)
    port map(
      ins => fork80_outs_1,
      ins_valid => fork80_outs_1_valid,
      ins_ready => fork80_outs_1_ready,
      clk => clk,
      rst => rst,
      outs => buffer225_outs,
      outs_valid => buffer225_outs_valid,
      outs_ready => buffer225_outs_ready
    );

  init132 : entity work.tehb_init(arch) generic map(32, 0)
    port map(
      ins => extsi43_outs,
      ins_valid => extsi43_outs_valid,
      ins_ready => extsi43_outs_ready,
      clk => clk,
      rst => rst,
      outs => init132_outs,
      outs_valid => init132_outs_valid,
      outs_ready => init132_outs_ready
    );

  buffer9 : entity work.tfifo_dataless(arch) generic map(1)
    port map(
      ins_valid => unbundle7_outs_0_valid,
      ins_ready => unbundle7_outs_0_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer9_outs_valid,
      outs_ready => buffer9_outs_ready
    );

  init133 : entity work.tehb_dataless_init(arch)
    port map(
      ins_valid => buffer9_outs_valid,
      ins_ready => buffer9_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => init133_outs_valid,
      outs_ready => init133_outs_ready
    );

  init134 : entity work.tehb_dataless_init(arch)
    port map(
      ins_valid => init133_outs_valid,
      ins_ready => init133_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => init134_outs_valid,
      outs_ready => init134_outs_ready
    );

  sink64 : entity work.sink_dataless(arch)
    port map(
      ins_valid => init134_outs_valid,
      ins_ready => init134_outs_ready,
      clk => clk,
      rst => rst
    );

  cond_br157 : entity work.cond_br_dataless(arch)
    port map(
      condition => buffer226_outs,
      condition_valid => buffer226_outs_valid,
      condition_ready => buffer226_outs_ready,
      data_valid => fork65_outs_0_valid,
      data_ready => fork65_outs_0_ready,
      clk => clk,
      rst => rst,
      trueOut_valid => cond_br157_trueOut_valid,
      trueOut_ready => cond_br157_trueOut_ready,
      falseOut_valid => cond_br157_falseOut_valid,
      falseOut_ready => cond_br157_falseOut_ready
    );

  buffer226 : entity work.tfifo(arch) generic map(1, 1)
    port map(
      ins => fork78_outs_1,
      ins_valid => fork78_outs_1_valid,
      ins_ready => fork78_outs_1_ready,
      clk => clk,
      rst => rst,
      outs => buffer226_outs,
      outs_valid => buffer226_outs_valid,
      outs_ready => buffer226_outs_ready
    );

  sink65 : entity work.sink_dataless(arch)
    port map(
      ins_valid => cond_br157_trueOut_valid,
      ins_ready => cond_br157_trueOut_ready,
      clk => clk,
      rst => rst
    );

  cond_br158 : entity work.cond_br_dataless(arch)
    port map(
      condition => buffer227_outs,
      condition_valid => buffer227_outs_valid,
      condition_ready => buffer227_outs_ready,
      data_valid => fork64_outs_0_valid,
      data_ready => fork64_outs_0_ready,
      clk => clk,
      rst => rst,
      trueOut_valid => cond_br158_trueOut_valid,
      trueOut_ready => cond_br158_trueOut_ready,
      falseOut_valid => cond_br158_falseOut_valid,
      falseOut_ready => cond_br158_falseOut_ready
    );

  buffer227 : entity work.tfifo(arch) generic map(1, 1)
    port map(
      ins => fork79_outs_1,
      ins_valid => fork79_outs_1_valid,
      ins_ready => fork79_outs_1_ready,
      clk => clk,
      rst => rst,
      outs => buffer227_outs,
      outs_valid => buffer227_outs_valid,
      outs_ready => buffer227_outs_ready
    );

  sink66 : entity work.sink_dataless(arch)
    port map(
      ins_valid => cond_br158_trueOut_valid,
      ins_ready => cond_br158_trueOut_ready,
      clk => clk,
      rst => rst
    );

  source15 : entity work.source(arch)
    port map(
      clk => clk,
      rst => rst,
      outs_valid => source15_outs_valid,
      outs_ready => source15_outs_ready
    );

  mux133 : entity work.mux_dataless(arch) generic map(2, 1)
    port map(
      index => buffer228_outs,
      index_valid => buffer228_outs_valid,
      index_ready => buffer228_outs_ready,
      ins_valid(0) => cond_br157_falseOut_valid,
      ins_valid(1) => source15_outs_valid,
      ins_ready(0) => cond_br157_falseOut_ready,
      ins_ready(1) => source15_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => mux133_outs_valid,
      outs_ready => mux133_outs_ready
    );

  buffer228 : entity work.tfifo(arch) generic map(1, 1)
    port map(
      ins => fork78_outs_0,
      ins_valid => fork78_outs_0_valid,
      ins_ready => fork78_outs_0_ready,
      clk => clk,
      rst => rst,
      outs => buffer228_outs,
      outs_valid => buffer228_outs_valid,
      outs_ready => buffer228_outs_ready
    );

  source16 : entity work.source(arch)
    port map(
      clk => clk,
      rst => rst,
      outs_valid => source16_outs_valid,
      outs_ready => source16_outs_ready
    );

  mux134 : entity work.mux_dataless(arch) generic map(2, 1)
    port map(
      index => buffer229_outs,
      index_valid => buffer229_outs_valid,
      index_ready => buffer229_outs_ready,
      ins_valid(0) => cond_br158_falseOut_valid,
      ins_valid(1) => source16_outs_valid,
      ins_ready(0) => cond_br158_falseOut_ready,
      ins_ready(1) => source16_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => mux134_outs_valid,
      outs_ready => mux134_outs_ready
    );

  buffer229 : entity work.tfifo(arch) generic map(1, 1)
    port map(
      ins => fork79_outs_0,
      ins_valid => fork79_outs_0_valid,
      ins_ready => fork79_outs_0_ready,
      clk => clk,
      rst => rst,
      outs => buffer229_outs,
      outs_valid => buffer229_outs_valid,
      outs_ready => buffer229_outs_ready
    );

  buffer103 : entity work.tehb_dataless(arch)
    port map(
      ins_valid => mux133_outs_valid,
      ins_ready => mux133_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer103_outs_valid,
      outs_ready => buffer103_outs_ready
    );

  buffer104 : entity work.tehb_dataless(arch)
    port map(
      ins_valid => mux134_outs_valid,
      ins_ready => mux134_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer104_outs_valid,
      outs_ready => buffer104_outs_ready
    );

  join4 : entity work.join_handshake(arch) generic map(2)
    port map(
      ins_valid(0) => buffer103_outs_valid,
      ins_valid(1) => buffer104_outs_valid,
      ins_ready(0) => buffer103_outs_ready,
      ins_ready(1) => buffer104_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => join4_outs_valid,
      outs_ready => join4_outs_ready
    );

  gate9 : entity work.gate(arch) generic map(2, 32)
    port map(
      ins(0) => buffer230_outs,
      ins_valid(0) => buffer230_outs_valid,
      ins_valid(1) => join4_outs_valid,
      ins_ready(0) => buffer230_outs_ready,
      ins_ready(1) => join4_outs_ready,
      clk => clk,
      rst => rst,
      outs => gate9_outs,
      outs_valid => gate9_outs_valid,
      outs_ready => gate9_outs_ready
    );

  buffer230 : entity work.tfifo(arch) generic map(1, 32)
    port map(
      ins => fork74_outs_1,
      ins_valid => fork74_outs_1_valid,
      ins_ready => fork74_outs_1_ready,
      clk => clk,
      rst => rst,
      outs => buffer230_outs,
      outs_valid => buffer230_outs_valid,
      outs_ready => buffer230_outs_ready
    );

  trunci5 : entity work.trunci(arch) generic map(32, 7)
    port map(
      ins => gate9_outs,
      ins_valid => gate9_outs_valid,
      ins_ready => gate9_outs_ready,
      clk => clk,
      rst => rst,
      outs => trunci5_outs,
      outs_valid => trunci5_outs_valid,
      outs_ready => trunci5_outs_ready
    );

  load3 : entity work.load(arch) generic map(32, 7)
    port map(
      addrIn => trunci5_outs,
      addrIn_valid => trunci5_outs_valid,
      addrIn_ready => trunci5_outs_ready,
      dataFromMem => mem_controller0_ldData_0,
      dataFromMem_valid => mem_controller0_ldData_0_valid,
      dataFromMem_ready => mem_controller0_ldData_0_ready,
      clk => clk,
      rst => rst,
      addrOut => load3_addrOut,
      addrOut_valid => load3_addrOut_valid,
      addrOut_ready => load3_addrOut_ready,
      dataOut => load3_dataOut,
      dataOut_valid => load3_dataOut_valid,
      dataOut_ready => load3_dataOut_ready
    );

  fork81 : entity work.handshake_fork(arch) generic map(2, 32)
    port map(
      ins => load3_dataOut,
      ins_valid => load3_dataOut_valid,
      ins_ready => load3_dataOut_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork81_outs_0,
      outs(1) => fork81_outs_1,
      outs_valid(0) => fork81_outs_0_valid,
      outs_valid(1) => fork81_outs_1_valid,
      outs_ready(0) => fork81_outs_0_ready,
      outs_ready(1) => fork81_outs_1_ready
    );

  gate10 : entity work.gate(arch) generic map(2, 32)
    port map(
      ins(0) => buffer231_outs,
      ins_valid(0) => buffer231_outs_valid,
      ins_valid(1) => fork61_outs_0_valid,
      ins_ready(0) => buffer231_outs_ready,
      ins_ready(1) => fork61_outs_0_ready,
      clk => clk,
      rst => rst,
      outs => gate10_outs,
      outs_valid => gate10_outs_valid,
      outs_ready => gate10_outs_ready
    );

  buffer231 : entity work.tfifo(arch) generic map(1, 32)
    port map(
      ins => fork74_outs_2,
      ins_valid => fork74_outs_2_valid,
      ins_ready => fork74_outs_2_ready,
      clk => clk,
      rst => rst,
      outs => buffer231_outs,
      outs_valid => buffer231_outs_valid,
      outs_ready => buffer231_outs_ready
    );

  fork82 : entity work.handshake_fork(arch) generic map(2, 32)
    port map(
      ins => gate10_outs,
      ins_valid => gate10_outs_valid,
      ins_ready => gate10_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork82_outs_0,
      outs(1) => fork82_outs_1,
      outs_valid(0) => fork82_outs_0_valid,
      outs_valid(1) => fork82_outs_1_valid,
      outs_ready(0) => fork82_outs_0_ready,
      outs_ready(1) => fork82_outs_1_ready
    );

  cmpi13 : entity work.handshake_cmpi_0(arch) generic map(32)
    port map(
      lhs => fork82_outs_1,
      lhs_valid => fork82_outs_1_valid,
      lhs_ready => fork82_outs_1_ready,
      rhs => extsi37_outs,
      rhs_valid => extsi37_outs_valid,
      rhs_ready => extsi37_outs_ready,
      clk => clk,
      rst => rst,
      result => cmpi13_result,
      result_valid => cmpi13_result_valid,
      result_ready => cmpi13_result_ready
    );

  fork83 : entity work.handshake_fork(arch) generic map(2, 1)
    port map(
      ins => cmpi13_result,
      ins_valid => cmpi13_result_valid,
      ins_ready => cmpi13_result_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork83_outs_0,
      outs(1) => fork83_outs_1,
      outs_valid(0) => fork83_outs_0_valid,
      outs_valid(1) => fork83_outs_1_valid,
      outs_ready(0) => fork83_outs_0_ready,
      outs_ready(1) => fork83_outs_1_ready
    );

  cmpi14 : entity work.handshake_cmpi_0(arch) generic map(32)
    port map(
      lhs => fork82_outs_0,
      lhs_valid => fork82_outs_0_valid,
      lhs_ready => fork82_outs_0_ready,
      rhs => buffer234_outs,
      rhs_valid => buffer234_outs_valid,
      rhs_ready => buffer234_outs_ready,
      clk => clk,
      rst => rst,
      result => cmpi14_result,
      result_valid => cmpi14_result_valid,
      result_ready => cmpi14_result_ready
    );

  buffer234 : entity work.tfifo(arch) generic map(1, 32)
    port map(
      ins => fork63_outs_0,
      ins_valid => fork63_outs_0_valid,
      ins_ready => fork63_outs_0_ready,
      clk => clk,
      rst => rst,
      outs => buffer234_outs,
      outs_valid => buffer234_outs_valid,
      outs_ready => buffer234_outs_ready
    );

  fork84 : entity work.handshake_fork(arch) generic map(2, 1)
    port map(
      ins => cmpi14_result,
      ins_valid => cmpi14_result_valid,
      ins_ready => cmpi14_result_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork84_outs_0,
      outs(1) => fork84_outs_1,
      outs_valid(0) => fork84_outs_0_valid,
      outs_valid(1) => fork84_outs_1_valid,
      outs_ready(0) => fork84_outs_0_ready,
      outs_ready(1) => fork84_outs_1_ready
    );

  gate11 : entity work.gate(arch) generic map(2, 32)
    port map(
      ins(0) => buffer235_outs,
      ins_valid(0) => buffer235_outs_valid,
      ins_valid(1) => fork68_outs_0_valid,
      ins_ready(0) => buffer235_outs_ready,
      ins_ready(1) => fork68_outs_0_ready,
      clk => clk,
      rst => rst,
      outs => gate11_outs,
      outs_valid => gate11_outs_valid,
      outs_ready => gate11_outs_ready
    );

  buffer235 : entity work.tfifo(arch) generic map(1, 32)
    port map(
      ins => fork74_outs_3,
      ins_valid => fork74_outs_3_valid,
      ins_ready => fork74_outs_3_ready,
      clk => clk,
      rst => rst,
      outs => buffer235_outs,
      outs_valid => buffer235_outs_valid,
      outs_ready => buffer235_outs_ready
    );

  fork85 : entity work.handshake_fork(arch) generic map(2, 32)
    port map(
      ins => gate11_outs,
      ins_valid => gate11_outs_valid,
      ins_ready => gate11_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork85_outs_0,
      outs(1) => fork85_outs_1,
      outs_valid(0) => fork85_outs_0_valid,
      outs_valid(1) => fork85_outs_1_valid,
      outs_ready(0) => fork85_outs_0_ready,
      outs_ready(1) => fork85_outs_1_ready
    );

  cmpi15 : entity work.handshake_cmpi_0(arch) generic map(32)
    port map(
      lhs => buffer236_outs,
      lhs_valid => buffer236_outs_valid,
      lhs_ready => buffer236_outs_ready,
      rhs => fork69_outs_0,
      rhs_valid => fork69_outs_0_valid,
      rhs_ready => fork69_outs_0_ready,
      clk => clk,
      rst => rst,
      result => cmpi15_result,
      result_valid => cmpi15_result_valid,
      result_ready => cmpi15_result_ready
    );

  buffer236 : entity work.tfifo(arch) generic map(1, 32)
    port map(
      ins => fork85_outs_1,
      ins_valid => fork85_outs_1_valid,
      ins_ready => fork85_outs_1_ready,
      clk => clk,
      rst => rst,
      outs => buffer236_outs,
      outs_valid => buffer236_outs_valid,
      outs_ready => buffer236_outs_ready
    );

  fork86 : entity work.handshake_fork(arch) generic map(2, 1)
    port map(
      ins => cmpi15_result,
      ins_valid => cmpi15_result_valid,
      ins_ready => cmpi15_result_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork86_outs_0,
      outs(1) => fork86_outs_1,
      outs_valid(0) => fork86_outs_0_valid,
      outs_valid(1) => fork86_outs_1_valid,
      outs_ready(0) => fork86_outs_0_ready,
      outs_ready(1) => fork86_outs_1_ready
    );

  cmpi16 : entity work.handshake_cmpi_0(arch) generic map(32)
    port map(
      lhs => buffer238_outs,
      lhs_valid => buffer238_outs_valid,
      lhs_ready => buffer238_outs_ready,
      rhs => fork70_outs_0,
      rhs_valid => fork70_outs_0_valid,
      rhs_ready => fork70_outs_0_ready,
      clk => clk,
      rst => rst,
      result => cmpi16_result,
      result_valid => cmpi16_result_valid,
      result_ready => cmpi16_result_ready
    );

  buffer238 : entity work.tfifo(arch) generic map(1, 32)
    port map(
      ins => fork85_outs_0,
      ins_valid => fork85_outs_0_valid,
      ins_ready => fork85_outs_0_ready,
      clk => clk,
      rst => rst,
      outs => buffer238_outs,
      outs_valid => buffer238_outs_valid,
      outs_ready => buffer238_outs_ready
    );

  fork87 : entity work.handshake_fork(arch) generic map(2, 1)
    port map(
      ins => cmpi16_result,
      ins_valid => cmpi16_result_valid,
      ins_ready => cmpi16_result_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork87_outs_0,
      outs(1) => fork87_outs_1,
      outs_valid(0) => fork87_outs_0_valid,
      outs_valid(1) => fork87_outs_1_valid,
      outs_ready(0) => fork87_outs_0_ready,
      outs_ready(1) => fork87_outs_1_ready
    );

  gate12 : entity work.gate(arch) generic map(2, 32)
    port map(
      ins(0) => buffer240_outs,
      ins_valid(0) => buffer240_outs_valid,
      ins_valid(1) => fork56_outs_0_valid,
      ins_ready(0) => buffer240_outs_ready,
      ins_ready(1) => fork56_outs_0_ready,
      clk => clk,
      rst => rst,
      outs => gate12_outs,
      outs_valid => gate12_outs_valid,
      outs_ready => gate12_outs_ready
    );

  buffer240 : entity work.tfifo(arch) generic map(1, 32)
    port map(
      ins => fork74_outs_4,
      ins_valid => fork74_outs_4_valid,
      ins_ready => fork74_outs_4_ready,
      clk => clk,
      rst => rst,
      outs => buffer240_outs,
      outs_valid => buffer240_outs_valid,
      outs_ready => buffer240_outs_ready
    );

  fork88 : entity work.handshake_fork(arch) generic map(2, 32)
    port map(
      ins => gate12_outs,
      ins_valid => gate12_outs_valid,
      ins_ready => gate12_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork88_outs_0,
      outs(1) => fork88_outs_1,
      outs_valid(0) => fork88_outs_0_valid,
      outs_valid(1) => fork88_outs_1_valid,
      outs_ready(0) => fork88_outs_0_ready,
      outs_ready(1) => fork88_outs_1_ready
    );

  cmpi17 : entity work.handshake_cmpi_0(arch) generic map(32)
    port map(
      lhs => fork88_outs_1,
      lhs_valid => fork88_outs_1_valid,
      lhs_ready => fork88_outs_1_ready,
      rhs => extsi36_outs,
      rhs_valid => extsi36_outs_valid,
      rhs_ready => extsi36_outs_ready,
      clk => clk,
      rst => rst,
      result => cmpi17_result,
      result_valid => cmpi17_result_valid,
      result_ready => cmpi17_result_ready
    );

  fork89 : entity work.handshake_fork(arch) generic map(2, 1)
    port map(
      ins => cmpi17_result,
      ins_valid => cmpi17_result_valid,
      ins_ready => cmpi17_result_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork89_outs_0,
      outs(1) => fork89_outs_1,
      outs_valid(0) => fork89_outs_0_valid,
      outs_valid(1) => fork89_outs_1_valid,
      outs_ready(0) => fork89_outs_0_ready,
      outs_ready(1) => fork89_outs_1_ready
    );

  cmpi18 : entity work.handshake_cmpi_0(arch) generic map(32)
    port map(
      lhs => fork88_outs_0,
      lhs_valid => fork88_outs_0_valid,
      lhs_ready => fork88_outs_0_ready,
      rhs => buffer243_outs,
      rhs_valid => buffer243_outs_valid,
      rhs_ready => buffer243_outs_ready,
      clk => clk,
      rst => rst,
      result => cmpi18_result,
      result_valid => cmpi18_result_valid,
      result_ready => cmpi18_result_ready
    );

  buffer243 : entity work.tfifo(arch) generic map(1, 32)
    port map(
      ins => fork55_outs_0,
      ins_valid => fork55_outs_0_valid,
      ins_ready => fork55_outs_0_ready,
      clk => clk,
      rst => rst,
      outs => buffer243_outs,
      outs_valid => buffer243_outs_valid,
      outs_ready => buffer243_outs_ready
    );

  fork90 : entity work.handshake_fork(arch) generic map(2, 1)
    port map(
      ins => cmpi18_result,
      ins_valid => cmpi18_result_valid,
      ins_ready => cmpi18_result_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork90_outs_0,
      outs(1) => fork90_outs_1,
      outs_valid(0) => fork90_outs_0_valid,
      outs_valid(1) => fork90_outs_1_valid,
      outs_ready(0) => fork90_outs_0_ready,
      outs_ready(1) => fork90_outs_1_ready
    );

  buffer10 : entity work.tfifo(arch) generic map(1, 8)
    port map(
      ins => fork73_outs_1,
      ins_valid => fork73_outs_1_valid,
      ins_ready => fork73_outs_1_ready,
      clk => clk,
      rst => rst,
      outs => buffer10_outs,
      outs_valid => buffer10_outs_valid,
      outs_ready => buffer10_outs_ready
    );

  fork91 : entity work.handshake_fork(arch) generic map(2, 8)
    port map(
      ins => buffer10_outs,
      ins_valid => buffer10_outs_valid,
      ins_ready => buffer10_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork91_outs_0,
      outs(1) => fork91_outs_1,
      outs_valid(0) => fork91_outs_0_valid,
      outs_valid(1) => fork91_outs_1_valid,
      outs_ready(0) => fork91_outs_0_ready,
      outs_ready(1) => fork91_outs_1_ready
    );

  extsi44 : entity work.extsi(arch) generic map(8, 32)
    port map(
      ins => buffer245_outs,
      ins_valid => buffer245_outs_valid,
      ins_ready => buffer245_outs_ready,
      clk => clk,
      rst => rst,
      outs => extsi44_outs,
      outs_valid => extsi44_outs_valid,
      outs_ready => extsi44_outs_ready
    );

  buffer245 : entity work.tfifo(arch) generic map(1, 8)
    port map(
      ins => fork91_outs_1,
      ins_valid => fork91_outs_1_valid,
      ins_ready => fork91_outs_1_ready,
      clk => clk,
      rst => rst,
      outs => buffer245_outs,
      outs_valid => buffer245_outs_valid,
      outs_ready => buffer245_outs_ready
    );

  init135 : entity work.tehb_init(arch) generic map(32, 0)
    port map(
      ins => extsi44_outs,
      ins_valid => extsi44_outs_valid,
      ins_ready => extsi44_outs_ready,
      clk => clk,
      rst => rst,
      outs => init135_outs,
      outs_valid => init135_outs_valid,
      outs_ready => init135_outs_ready
    );

  buffer11 : entity work.tfifo_dataless(arch) generic map(1)
    port map(
      ins_valid => store1_doneOut_valid,
      ins_ready => store1_doneOut_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer11_outs_valid,
      outs_ready => buffer11_outs_ready
    );

  init136 : entity work.tehb_dataless_init(arch)
    port map(
      ins_valid => buffer11_outs_valid,
      ins_ready => buffer11_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => init136_outs_valid,
      outs_ready => init136_outs_ready
    );

  fork92 : entity work.fork_dataless(arch) generic map(2)
    port map(
      ins_valid => init136_outs_valid,
      ins_ready => init136_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid(0) => fork92_outs_0_valid,
      outs_valid(1) => fork92_outs_1_valid,
      outs_ready(0) => fork92_outs_0_ready,
      outs_ready(1) => fork92_outs_1_ready
    );

  init137 : entity work.tehb_dataless_init(arch)
    port map(
      ins_valid => fork92_outs_0_valid,
      ins_ready => fork92_outs_0_ready,
      clk => clk,
      rst => rst,
      outs_valid => init137_outs_valid,
      outs_ready => init137_outs_ready
    );

  sink67 : entity work.sink_dataless(arch)
    port map(
      ins_valid => init137_outs_valid,
      ins_ready => init137_outs_ready,
      clk => clk,
      rst => rst
    );

  cond_br159 : entity work.cond_br_dataless(arch)
    port map(
      condition => fork83_outs_1,
      condition_valid => fork83_outs_1_valid,
      condition_ready => fork83_outs_1_ready,
      data_valid => fork67_outs_0_valid,
      data_ready => fork67_outs_0_ready,
      clk => clk,
      rst => rst,
      trueOut_valid => cond_br159_trueOut_valid,
      trueOut_ready => cond_br159_trueOut_ready,
      falseOut_valid => cond_br159_falseOut_valid,
      falseOut_ready => cond_br159_falseOut_ready
    );

  sink68 : entity work.sink_dataless(arch)
    port map(
      ins_valid => cond_br159_trueOut_valid,
      ins_ready => cond_br159_trueOut_ready,
      clk => clk,
      rst => rst
    );

  cond_br160 : entity work.cond_br_dataless(arch)
    port map(
      condition => buffer247_outs,
      condition_valid => buffer247_outs_valid,
      condition_ready => buffer247_outs_ready,
      data_valid => fork66_outs_0_valid,
      data_ready => fork66_outs_0_ready,
      clk => clk,
      rst => rst,
      trueOut_valid => cond_br160_trueOut_valid,
      trueOut_ready => cond_br160_trueOut_ready,
      falseOut_valid => cond_br160_falseOut_valid,
      falseOut_ready => cond_br160_falseOut_ready
    );

  buffer247 : entity work.tfifo(arch) generic map(1, 1)
    port map(
      ins => fork84_outs_1,
      ins_valid => fork84_outs_1_valid,
      ins_ready => fork84_outs_1_ready,
      clk => clk,
      rst => rst,
      outs => buffer247_outs,
      outs_valid => buffer247_outs_valid,
      outs_ready => buffer247_outs_ready
    );

  sink69 : entity work.sink_dataless(arch)
    port map(
      ins_valid => cond_br160_trueOut_valid,
      ins_ready => cond_br160_trueOut_ready,
      clk => clk,
      rst => rst
    );

  source17 : entity work.source(arch)
    port map(
      clk => clk,
      rst => rst,
      outs_valid => source17_outs_valid,
      outs_ready => source17_outs_ready
    );

  mux135 : entity work.mux_dataless(arch) generic map(2, 1)
    port map(
      index => buffer248_outs,
      index_valid => buffer248_outs_valid,
      index_ready => buffer248_outs_ready,
      ins_valid(0) => cond_br159_falseOut_valid,
      ins_valid(1) => source17_outs_valid,
      ins_ready(0) => cond_br159_falseOut_ready,
      ins_ready(1) => source17_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => mux135_outs_valid,
      outs_ready => mux135_outs_ready
    );

  buffer248 : entity work.tfifo(arch) generic map(1, 1)
    port map(
      ins => fork83_outs_0,
      ins_valid => fork83_outs_0_valid,
      ins_ready => fork83_outs_0_ready,
      clk => clk,
      rst => rst,
      outs => buffer248_outs,
      outs_valid => buffer248_outs_valid,
      outs_ready => buffer248_outs_ready
    );

  source18 : entity work.source(arch)
    port map(
      clk => clk,
      rst => rst,
      outs_valid => source18_outs_valid,
      outs_ready => source18_outs_ready
    );

  mux136 : entity work.mux_dataless(arch) generic map(2, 1)
    port map(
      index => buffer249_outs,
      index_valid => buffer249_outs_valid,
      index_ready => buffer249_outs_ready,
      ins_valid(0) => cond_br160_falseOut_valid,
      ins_valid(1) => source18_outs_valid,
      ins_ready(0) => cond_br160_falseOut_ready,
      ins_ready(1) => source18_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => mux136_outs_valid,
      outs_ready => mux136_outs_ready
    );

  buffer249 : entity work.tfifo(arch) generic map(1, 1)
    port map(
      ins => fork84_outs_0,
      ins_valid => fork84_outs_0_valid,
      ins_ready => fork84_outs_0_ready,
      clk => clk,
      rst => rst,
      outs => buffer249_outs,
      outs_valid => buffer249_outs_valid,
      outs_ready => buffer249_outs_ready
    );

  buffer105 : entity work.tehb_dataless(arch)
    port map(
      ins_valid => mux135_outs_valid,
      ins_ready => mux135_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer105_outs_valid,
      outs_ready => buffer105_outs_ready
    );

  buffer106 : entity work.tehb_dataless(arch)
    port map(
      ins_valid => mux136_outs_valid,
      ins_ready => mux136_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer106_outs_valid,
      outs_ready => buffer106_outs_ready
    );

  join5 : entity work.join_handshake(arch) generic map(2)
    port map(
      ins_valid(0) => buffer105_outs_valid,
      ins_valid(1) => buffer106_outs_valid,
      ins_ready(0) => buffer105_outs_ready,
      ins_ready(1) => buffer106_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => join5_outs_valid,
      outs_ready => join5_outs_ready
    );

  cond_br161 : entity work.cond_br_dataless(arch)
    port map(
      condition => buffer250_outs,
      condition_valid => buffer250_outs_valid,
      condition_ready => buffer250_outs_ready,
      data_valid => fork72_outs_0_valid,
      data_ready => fork72_outs_0_ready,
      clk => clk,
      rst => rst,
      trueOut_valid => cond_br161_trueOut_valid,
      trueOut_ready => cond_br161_trueOut_ready,
      falseOut_valid => cond_br161_falseOut_valid,
      falseOut_ready => cond_br161_falseOut_ready
    );

  buffer250 : entity work.tfifo(arch) generic map(1, 1)
    port map(
      ins => fork86_outs_1,
      ins_valid => fork86_outs_1_valid,
      ins_ready => fork86_outs_1_ready,
      clk => clk,
      rst => rst,
      outs => buffer250_outs,
      outs_valid => buffer250_outs_valid,
      outs_ready => buffer250_outs_ready
    );

  sink70 : entity work.sink_dataless(arch)
    port map(
      ins_valid => cond_br161_trueOut_valid,
      ins_ready => cond_br161_trueOut_ready,
      clk => clk,
      rst => rst
    );

  cond_br162 : entity work.cond_br_dataless(arch)
    port map(
      condition => buffer251_outs,
      condition_valid => buffer251_outs_valid,
      condition_ready => buffer251_outs_ready,
      data_valid => fork71_outs_0_valid,
      data_ready => fork71_outs_0_ready,
      clk => clk,
      rst => rst,
      trueOut_valid => cond_br162_trueOut_valid,
      trueOut_ready => cond_br162_trueOut_ready,
      falseOut_valid => cond_br162_falseOut_valid,
      falseOut_ready => cond_br162_falseOut_ready
    );

  buffer251 : entity work.tfifo(arch) generic map(1, 1)
    port map(
      ins => fork87_outs_1,
      ins_valid => fork87_outs_1_valid,
      ins_ready => fork87_outs_1_ready,
      clk => clk,
      rst => rst,
      outs => buffer251_outs,
      outs_valid => buffer251_outs_valid,
      outs_ready => buffer251_outs_ready
    );

  sink71 : entity work.sink_dataless(arch)
    port map(
      ins_valid => cond_br162_trueOut_valid,
      ins_ready => cond_br162_trueOut_ready,
      clk => clk,
      rst => rst
    );

  source19 : entity work.source(arch)
    port map(
      clk => clk,
      rst => rst,
      outs_valid => source19_outs_valid,
      outs_ready => source19_outs_ready
    );

  mux137 : entity work.mux_dataless(arch) generic map(2, 1)
    port map(
      index => buffer252_outs,
      index_valid => buffer252_outs_valid,
      index_ready => buffer252_outs_ready,
      ins_valid(0) => cond_br161_falseOut_valid,
      ins_valid(1) => source19_outs_valid,
      ins_ready(0) => cond_br161_falseOut_ready,
      ins_ready(1) => source19_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => mux137_outs_valid,
      outs_ready => mux137_outs_ready
    );

  buffer252 : entity work.tfifo(arch) generic map(1, 1)
    port map(
      ins => fork86_outs_0,
      ins_valid => fork86_outs_0_valid,
      ins_ready => fork86_outs_0_ready,
      clk => clk,
      rst => rst,
      outs => buffer252_outs,
      outs_valid => buffer252_outs_valid,
      outs_ready => buffer252_outs_ready
    );

  source20 : entity work.source(arch)
    port map(
      clk => clk,
      rst => rst,
      outs_valid => source20_outs_valid,
      outs_ready => source20_outs_ready
    );

  mux138 : entity work.mux_dataless(arch) generic map(2, 1)
    port map(
      index => buffer253_outs,
      index_valid => buffer253_outs_valid,
      index_ready => buffer253_outs_ready,
      ins_valid(0) => cond_br162_falseOut_valid,
      ins_valid(1) => source20_outs_valid,
      ins_ready(0) => cond_br162_falseOut_ready,
      ins_ready(1) => source20_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => mux138_outs_valid,
      outs_ready => mux138_outs_ready
    );

  buffer253 : entity work.tfifo(arch) generic map(1, 1)
    port map(
      ins => fork87_outs_0,
      ins_valid => fork87_outs_0_valid,
      ins_ready => fork87_outs_0_ready,
      clk => clk,
      rst => rst,
      outs => buffer253_outs,
      outs_valid => buffer253_outs_valid,
      outs_ready => buffer253_outs_ready
    );

  buffer107 : entity work.tehb_dataless(arch)
    port map(
      ins_valid => mux137_outs_valid,
      ins_ready => mux137_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer107_outs_valid,
      outs_ready => buffer107_outs_ready
    );

  buffer108 : entity work.tehb_dataless(arch)
    port map(
      ins_valid => mux138_outs_valid,
      ins_ready => mux138_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer108_outs_valid,
      outs_ready => buffer108_outs_ready
    );

  join6 : entity work.join_handshake(arch) generic map(2)
    port map(
      ins_valid(0) => buffer107_outs_valid,
      ins_valid(1) => buffer108_outs_valid,
      ins_ready(0) => buffer107_outs_ready,
      ins_ready(1) => buffer108_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => join6_outs_valid,
      outs_ready => join6_outs_ready
    );

  cond_br163 : entity work.cond_br_dataless(arch)
    port map(
      condition => buffer254_outs,
      condition_valid => buffer254_outs_valid,
      condition_ready => buffer254_outs_ready,
      data_valid => fork54_outs_0_valid,
      data_ready => fork54_outs_0_ready,
      clk => clk,
      rst => rst,
      trueOut_valid => cond_br163_trueOut_valid,
      trueOut_ready => cond_br163_trueOut_ready,
      falseOut_valid => cond_br163_falseOut_valid,
      falseOut_ready => cond_br163_falseOut_ready
    );

  buffer254 : entity work.tfifo(arch) generic map(1, 1)
    port map(
      ins => fork89_outs_1,
      ins_valid => fork89_outs_1_valid,
      ins_ready => fork89_outs_1_ready,
      clk => clk,
      rst => rst,
      outs => buffer254_outs,
      outs_valid => buffer254_outs_valid,
      outs_ready => buffer254_outs_ready
    );

  sink72 : entity work.sink_dataless(arch)
    port map(
      ins_valid => cond_br163_trueOut_valid,
      ins_ready => cond_br163_trueOut_ready,
      clk => clk,
      rst => rst
    );

  cond_br164 : entity work.cond_br_dataless(arch)
    port map(
      condition => buffer255_outs,
      condition_valid => buffer255_outs_valid,
      condition_ready => buffer255_outs_ready,
      data_valid => fork60_outs_0_valid,
      data_ready => fork60_outs_0_ready,
      clk => clk,
      rst => rst,
      trueOut_valid => cond_br164_trueOut_valid,
      trueOut_ready => cond_br164_trueOut_ready,
      falseOut_valid => cond_br164_falseOut_valid,
      falseOut_ready => cond_br164_falseOut_ready
    );

  buffer255 : entity work.tfifo(arch) generic map(1, 1)
    port map(
      ins => fork90_outs_1,
      ins_valid => fork90_outs_1_valid,
      ins_ready => fork90_outs_1_ready,
      clk => clk,
      rst => rst,
      outs => buffer255_outs,
      outs_valid => buffer255_outs_valid,
      outs_ready => buffer255_outs_ready
    );

  sink73 : entity work.sink_dataless(arch)
    port map(
      ins_valid => cond_br164_trueOut_valid,
      ins_ready => cond_br164_trueOut_ready,
      clk => clk,
      rst => rst
    );

  source21 : entity work.source(arch)
    port map(
      clk => clk,
      rst => rst,
      outs_valid => source21_outs_valid,
      outs_ready => source21_outs_ready
    );

  mux139 : entity work.mux_dataless(arch) generic map(2, 1)
    port map(
      index => buffer256_outs,
      index_valid => buffer256_outs_valid,
      index_ready => buffer256_outs_ready,
      ins_valid(0) => cond_br163_falseOut_valid,
      ins_valid(1) => source21_outs_valid,
      ins_ready(0) => cond_br163_falseOut_ready,
      ins_ready(1) => source21_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => mux139_outs_valid,
      outs_ready => mux139_outs_ready
    );

  buffer256 : entity work.tfifo(arch) generic map(1, 1)
    port map(
      ins => fork89_outs_0,
      ins_valid => fork89_outs_0_valid,
      ins_ready => fork89_outs_0_ready,
      clk => clk,
      rst => rst,
      outs => buffer256_outs,
      outs_valid => buffer256_outs_valid,
      outs_ready => buffer256_outs_ready
    );

  source22 : entity work.source(arch)
    port map(
      clk => clk,
      rst => rst,
      outs_valid => source22_outs_valid,
      outs_ready => source22_outs_ready
    );

  mux140 : entity work.mux_dataless(arch) generic map(2, 1)
    port map(
      index => buffer257_outs,
      index_valid => buffer257_outs_valid,
      index_ready => buffer257_outs_ready,
      ins_valid(0) => cond_br164_falseOut_valid,
      ins_valid(1) => source22_outs_valid,
      ins_ready(0) => cond_br164_falseOut_ready,
      ins_ready(1) => source22_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => mux140_outs_valid,
      outs_ready => mux140_outs_ready
    );

  buffer257 : entity work.tfifo(arch) generic map(1, 1)
    port map(
      ins => fork90_outs_0,
      ins_valid => fork90_outs_0_valid,
      ins_ready => fork90_outs_0_ready,
      clk => clk,
      rst => rst,
      outs => buffer257_outs,
      outs_valid => buffer257_outs_valid,
      outs_ready => buffer257_outs_ready
    );

  buffer109 : entity work.tehb_dataless(arch)
    port map(
      ins_valid => mux139_outs_valid,
      ins_ready => mux139_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer109_outs_valid,
      outs_ready => buffer109_outs_ready
    );

  buffer110 : entity work.tehb_dataless(arch)
    port map(
      ins_valid => mux140_outs_valid,
      ins_ready => mux140_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer110_outs_valid,
      outs_ready => buffer110_outs_ready
    );

  join7 : entity work.join_handshake(arch) generic map(2)
    port map(
      ins_valid(0) => buffer109_outs_valid,
      ins_valid(1) => buffer110_outs_valid,
      ins_ready(0) => buffer109_outs_ready,
      ins_ready(1) => buffer110_outs_ready,
      clk => clk,
      rst => rst,
      outs_valid => join7_outs_valid,
      outs_ready => join7_outs_ready
    );

  gate13 : entity work.gate(arch) generic map(4, 32)
    port map(
      ins(0) => buffer258_outs,
      ins_valid(0) => buffer258_outs_valid,
      ins_valid(1) => join5_outs_valid,
      ins_valid(2) => join6_outs_valid,
      ins_valid(3) => join7_outs_valid,
      ins_ready(0) => buffer258_outs_ready,
      ins_ready(1) => join5_outs_ready,
      ins_ready(2) => join6_outs_ready,
      ins_ready(3) => join7_outs_ready,
      clk => clk,
      rst => rst,
      outs => gate13_outs,
      outs_valid => gate13_outs_valid,
      outs_ready => gate13_outs_ready
    );

  buffer258 : entity work.tfifo(arch) generic map(1, 32)
    port map(
      ins => fork74_outs_5,
      ins_valid => fork74_outs_5_valid,
      ins_ready => fork74_outs_5_ready,
      clk => clk,
      rst => rst,
      outs => buffer258_outs,
      outs_valid => buffer258_outs_valid,
      outs_ready => buffer258_outs_ready
    );

  buffer111 : entity work.oehb(arch) generic map(32)
    port map(
      ins => gate13_outs,
      ins_valid => gate13_outs_valid,
      ins_ready => gate13_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer111_outs,
      outs_valid => buffer111_outs_valid,
      outs_ready => buffer111_outs_ready
    );

  trunci6 : entity work.trunci(arch) generic map(32, 7)
    port map(
      ins => buffer111_outs,
      ins_valid => buffer111_outs_valid,
      ins_ready => buffer111_outs_ready,
      clk => clk,
      rst => rst,
      outs => trunci6_outs,
      outs_valid => trunci6_outs_valid,
      outs_ready => trunci6_outs_ready
    );

  store1 : entity work.store(arch) generic map(32, 7)
    port map(
      addrIn => trunci6_outs,
      addrIn_valid => trunci6_outs_valid,
      addrIn_ready => trunci6_outs_ready,
      dataIn => fork81_outs_0,
      dataIn_valid => fork81_outs_0_valid,
      dataIn_ready => fork81_outs_0_ready,
      doneFromMem_valid => mem_controller1_stDone_0_valid,
      doneFromMem_ready => mem_controller1_stDone_0_ready,
      clk => clk,
      rst => rst,
      addrOut => store1_addrOut,
      addrOut_valid => store1_addrOut_valid,
      addrOut_ready => store1_addrOut_ready,
      dataToMem => store1_dataToMem,
      dataToMem_valid => store1_dataToMem_valid,
      dataToMem_ready => store1_dataToMem_ready,
      doneOut_valid => store1_doneOut_valid,
      doneOut_ready => store1_doneOut_ready
    );

  addi5 : entity work.addi(arch) generic map(9)
    port map(
      lhs => extsi39_outs,
      lhs_valid => extsi39_outs_valid,
      lhs_ready => extsi39_outs_ready,
      rhs => extsi42_outs,
      rhs_valid => extsi42_outs_valid,
      rhs_ready => extsi42_outs_ready,
      clk => clk,
      rst => rst,
      result => addi5_result,
      result_valid => addi5_result_valid,
      result_ready => addi5_result_ready
    );

  buffer112 : entity work.oehb(arch) generic map(9)
    port map(
      ins => addi5_result,
      ins_valid => addi5_result_valid,
      ins_ready => addi5_result_ready,
      clk => clk,
      rst => rst,
      outs => buffer112_outs,
      outs_valid => buffer112_outs_valid,
      outs_ready => buffer112_outs_ready
    );

  fork93 : entity work.handshake_fork(arch) generic map(2, 9)
    port map(
      ins => buffer112_outs,
      ins_valid => buffer112_outs_valid,
      ins_ready => buffer112_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork93_outs_0,
      outs(1) => fork93_outs_1,
      outs_valid(0) => fork93_outs_0_valid,
      outs_valid(1) => fork93_outs_1_valid,
      outs_ready(0) => fork93_outs_0_ready,
      outs_ready(1) => fork93_outs_1_ready
    );

  trunci7 : entity work.trunci(arch) generic map(9, 8)
    port map(
      ins => buffer260_outs,
      ins_valid => buffer260_outs_valid,
      ins_ready => buffer260_outs_ready,
      clk => clk,
      rst => rst,
      outs => trunci7_outs,
      outs_valid => trunci7_outs_valid,
      outs_ready => trunci7_outs_ready
    );

  buffer260 : entity work.tfifo(arch) generic map(1, 9)
    port map(
      ins => fork93_outs_0,
      ins_valid => fork93_outs_0_valid,
      ins_ready => fork93_outs_0_ready,
      clk => clk,
      rst => rst,
      outs => buffer260_outs,
      outs_valid => buffer260_outs_valid,
      outs_ready => buffer260_outs_ready
    );

  cmpi1 : entity work.handshake_cmpi_1(arch) generic map(9)
    port map(
      lhs => buffer261_outs,
      lhs_valid => buffer261_outs_valid,
      lhs_ready => buffer261_outs_ready,
      rhs => extsi41_outs,
      rhs_valid => extsi41_outs_valid,
      rhs_ready => extsi41_outs_ready,
      clk => clk,
      rst => rst,
      result => cmpi1_result,
      result_valid => cmpi1_result_valid,
      result_ready => cmpi1_result_ready
    );

  buffer261 : entity work.tfifo(arch) generic map(1, 9)
    port map(
      ins => fork93_outs_1,
      ins_valid => fork93_outs_1_valid,
      ins_ready => fork93_outs_1_ready,
      clk => clk,
      rst => rst,
      outs => buffer261_outs,
      outs_valid => buffer261_outs_valid,
      outs_ready => buffer261_outs_ready
    );

  buffer113 : entity work.oehb(arch) generic map(1)
    port map(
      ins => cmpi1_result,
      ins_valid => cmpi1_result_valid,
      ins_ready => cmpi1_result_ready,
      clk => clk,
      rst => rst,
      outs => buffer113_outs,
      outs_valid => buffer113_outs_valid,
      outs_ready => buffer113_outs_ready
    );

  fork94 : entity work.handshake_fork(arch) generic map(29, 1)
    port map(
      ins => buffer113_outs,
      ins_valid => buffer113_outs_valid,
      ins_ready => buffer113_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork94_outs_0,
      outs(1) => fork94_outs_1,
      outs(2) => fork94_outs_2,
      outs(3) => fork94_outs_3,
      outs(4) => fork94_outs_4,
      outs(5) => fork94_outs_5,
      outs(6) => fork94_outs_6,
      outs(7) => fork94_outs_7,
      outs(8) => fork94_outs_8,
      outs(9) => fork94_outs_9,
      outs(10) => fork94_outs_10,
      outs(11) => fork94_outs_11,
      outs(12) => fork94_outs_12,
      outs(13) => fork94_outs_13,
      outs(14) => fork94_outs_14,
      outs(15) => fork94_outs_15,
      outs(16) => fork94_outs_16,
      outs(17) => fork94_outs_17,
      outs(18) => fork94_outs_18,
      outs(19) => fork94_outs_19,
      outs(20) => fork94_outs_20,
      outs(21) => fork94_outs_21,
      outs(22) => fork94_outs_22,
      outs(23) => fork94_outs_23,
      outs(24) => fork94_outs_24,
      outs(25) => fork94_outs_25,
      outs(26) => fork94_outs_26,
      outs(27) => fork94_outs_27,
      outs(28) => fork94_outs_28,
      outs_valid(0) => fork94_outs_0_valid,
      outs_valid(1) => fork94_outs_1_valid,
      outs_valid(2) => fork94_outs_2_valid,
      outs_valid(3) => fork94_outs_3_valid,
      outs_valid(4) => fork94_outs_4_valid,
      outs_valid(5) => fork94_outs_5_valid,
      outs_valid(6) => fork94_outs_6_valid,
      outs_valid(7) => fork94_outs_7_valid,
      outs_valid(8) => fork94_outs_8_valid,
      outs_valid(9) => fork94_outs_9_valid,
      outs_valid(10) => fork94_outs_10_valid,
      outs_valid(11) => fork94_outs_11_valid,
      outs_valid(12) => fork94_outs_12_valid,
      outs_valid(13) => fork94_outs_13_valid,
      outs_valid(14) => fork94_outs_14_valid,
      outs_valid(15) => fork94_outs_15_valid,
      outs_valid(16) => fork94_outs_16_valid,
      outs_valid(17) => fork94_outs_17_valid,
      outs_valid(18) => fork94_outs_18_valid,
      outs_valid(19) => fork94_outs_19_valid,
      outs_valid(20) => fork94_outs_20_valid,
      outs_valid(21) => fork94_outs_21_valid,
      outs_valid(22) => fork94_outs_22_valid,
      outs_valid(23) => fork94_outs_23_valid,
      outs_valid(24) => fork94_outs_24_valid,
      outs_valid(25) => fork94_outs_25_valid,
      outs_valid(26) => fork94_outs_26_valid,
      outs_valid(27) => fork94_outs_27_valid,
      outs_valid(28) => fork94_outs_28_valid,
      outs_ready(0) => fork94_outs_0_ready,
      outs_ready(1) => fork94_outs_1_ready,
      outs_ready(2) => fork94_outs_2_ready,
      outs_ready(3) => fork94_outs_3_ready,
      outs_ready(4) => fork94_outs_4_ready,
      outs_ready(5) => fork94_outs_5_ready,
      outs_ready(6) => fork94_outs_6_ready,
      outs_ready(7) => fork94_outs_7_ready,
      outs_ready(8) => fork94_outs_8_ready,
      outs_ready(9) => fork94_outs_9_ready,
      outs_ready(10) => fork94_outs_10_ready,
      outs_ready(11) => fork94_outs_11_ready,
      outs_ready(12) => fork94_outs_12_ready,
      outs_ready(13) => fork94_outs_13_ready,
      outs_ready(14) => fork94_outs_14_ready,
      outs_ready(15) => fork94_outs_15_ready,
      outs_ready(16) => fork94_outs_16_ready,
      outs_ready(17) => fork94_outs_17_ready,
      outs_ready(18) => fork94_outs_18_ready,
      outs_ready(19) => fork94_outs_19_ready,
      outs_ready(20) => fork94_outs_20_ready,
      outs_ready(21) => fork94_outs_21_ready,
      outs_ready(22) => fork94_outs_22_ready,
      outs_ready(23) => fork94_outs_23_ready,
      outs_ready(24) => fork94_outs_24_ready,
      outs_ready(25) => fork94_outs_25_ready,
      outs_ready(26) => fork94_outs_26_ready,
      outs_ready(27) => fork94_outs_27_ready,
      outs_ready(28) => fork94_outs_28_ready
    );

  cond_br7 : entity work.cond_br(arch) generic map(8)
    port map(
      condition => fork94_outs_0,
      condition_valid => fork94_outs_0_valid,
      condition_ready => fork94_outs_0_ready,
      data => trunci7_outs,
      data_valid => trunci7_outs_valid,
      data_ready => trunci7_outs_ready,
      clk => clk,
      rst => rst,
      trueOut => cond_br7_trueOut,
      trueOut_valid => cond_br7_trueOut_valid,
      trueOut_ready => cond_br7_trueOut_ready,
      falseOut => cond_br7_falseOut,
      falseOut_valid => cond_br7_falseOut_valid,
      falseOut_ready => cond_br7_falseOut_ready
    );

  sink74 : entity work.sink(arch) generic map(8)
    port map(
      ins => cond_br7_falseOut,
      ins_valid => cond_br7_falseOut_valid,
      ins_ready => cond_br7_falseOut_ready,
      clk => clk,
      rst => rst
    );

  buffer100 : entity work.oehb(arch) generic map(3)
    port map(
      ins => mux4_outs,
      ins_valid => mux4_outs_valid,
      ins_ready => mux4_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer100_outs,
      outs_valid => buffer100_outs_valid,
      outs_ready => buffer100_outs_ready
    );

  buffer101 : entity work.tehb(arch) generic map(3)
    port map(
      ins => buffer100_outs,
      ins_valid => buffer100_outs_valid,
      ins_ready => buffer100_outs_ready,
      clk => clk,
      rst => rst,
      outs => buffer101_outs,
      outs_valid => buffer101_outs_valid,
      outs_ready => buffer101_outs_ready
    );

  cond_br8 : entity work.cond_br(arch) generic map(3)
    port map(
      condition => fork94_outs_1,
      condition_valid => fork94_outs_1_valid,
      condition_ready => fork94_outs_1_ready,
      data => buffer101_outs,
      data_valid => buffer101_outs_valid,
      data_ready => buffer101_outs_ready,
      clk => clk,
      rst => rst,
      trueOut => cond_br8_trueOut,
      trueOut_valid => cond_br8_trueOut_valid,
      trueOut_ready => cond_br8_trueOut_ready,
      falseOut => cond_br8_falseOut,
      falseOut_valid => cond_br8_falseOut_valid,
      falseOut_ready => cond_br8_falseOut_ready
    );

  buffer102 : entity work.oehb_dataless(arch)
    port map(
      ins_valid => fork76_outs_1_valid,
      ins_ready => fork76_outs_1_ready,
      clk => clk,
      rst => rst,
      outs_valid => buffer102_outs_valid,
      outs_ready => buffer102_outs_ready
    );

  cond_br9 : entity work.cond_br_dataless(arch)
    port map(
      condition => buffer264_outs,
      condition_valid => buffer264_outs_valid,
      condition_ready => buffer264_outs_ready,
      data_valid => buffer102_outs_valid,
      data_ready => buffer102_outs_ready,
      clk => clk,
      rst => rst,
      trueOut_valid => cond_br9_trueOut_valid,
      trueOut_ready => cond_br9_trueOut_ready,
      falseOut_valid => cond_br9_falseOut_valid,
      falseOut_ready => cond_br9_falseOut_ready
    );

  buffer264 : entity work.tfifo(arch) generic map(1, 1)
    port map(
      ins => fork94_outs_28,
      ins_valid => fork94_outs_28_valid,
      ins_ready => fork94_outs_28_ready,
      clk => clk,
      rst => rst,
      outs => buffer264_outs,
      outs_valid => buffer264_outs_valid,
      outs_ready => buffer264_outs_ready
    );

  cond_br259 : entity work.cond_br(arch) generic map(32)
    port map(
      condition => fork98_outs_3,
      condition_valid => fork98_outs_3_valid,
      condition_ready => fork98_outs_3_ready,
      data => cond_br244_falseOut,
      data_valid => cond_br244_falseOut_valid,
      data_ready => cond_br244_falseOut_ready,
      clk => clk,
      rst => rst,
      trueOut => cond_br259_trueOut,
      trueOut_valid => cond_br259_trueOut_valid,
      trueOut_ready => cond_br259_trueOut_ready,
      falseOut => cond_br259_falseOut,
      falseOut_valid => cond_br259_falseOut_valid,
      falseOut_ready => cond_br259_falseOut_ready
    );

  sink75 : entity work.sink(arch) generic map(32)
    port map(
      ins => cond_br259_falseOut,
      ins_valid => cond_br259_falseOut_valid,
      ins_ready => cond_br259_falseOut_ready,
      clk => clk,
      rst => rst
    );

  fork95 : entity work.handshake_fork(arch) generic map(3, 32)
    port map(
      ins => cond_br259_trueOut,
      ins_valid => cond_br259_trueOut_valid,
      ins_ready => cond_br259_trueOut_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork95_outs_0,
      outs(1) => fork95_outs_1,
      outs(2) => fork95_outs_2,
      outs_valid(0) => fork95_outs_0_valid,
      outs_valid(1) => fork95_outs_1_valid,
      outs_valid(2) => fork95_outs_2_valid,
      outs_ready(0) => fork95_outs_0_ready,
      outs_ready(1) => fork95_outs_1_ready,
      outs_ready(2) => fork95_outs_2_ready
    );

  cond_br260 : entity work.cond_br(arch) generic map(8)
    port map(
      condition => fork98_outs_7,
      condition_valid => fork98_outs_7_valid,
      condition_ready => fork98_outs_7_ready,
      data => cond_br246_falseOut,
      data_valid => cond_br246_falseOut_valid,
      data_ready => cond_br246_falseOut_ready,
      clk => clk,
      rst => rst,
      trueOut => cond_br260_trueOut,
      trueOut_valid => cond_br260_trueOut_valid,
      trueOut_ready => cond_br260_trueOut_ready,
      falseOut => cond_br260_falseOut,
      falseOut_valid => cond_br260_falseOut_valid,
      falseOut_ready => cond_br260_falseOut_ready
    );

  sink76 : entity work.sink(arch) generic map(8)
    port map(
      ins => cond_br260_falseOut,
      ins_valid => cond_br260_falseOut_valid,
      ins_ready => cond_br260_falseOut_ready,
      clk => clk,
      rst => rst
    );

  fork96 : entity work.handshake_fork(arch) generic map(3, 8)
    port map(
      ins => cond_br260_trueOut,
      ins_valid => cond_br260_trueOut_valid,
      ins_ready => cond_br260_trueOut_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork96_outs_0,
      outs(1) => fork96_outs_1,
      outs(2) => fork96_outs_2,
      outs_valid(0) => fork96_outs_0_valid,
      outs_valid(1) => fork96_outs_1_valid,
      outs_valid(2) => fork96_outs_2_valid,
      outs_ready(0) => fork96_outs_0_ready,
      outs_ready(1) => fork96_outs_1_ready,
      outs_ready(2) => fork96_outs_2_ready
    );

  extsi45 : entity work.extsi(arch) generic map(8, 11)
    port map(
      ins => fork96_outs_0,
      ins_valid => fork96_outs_0_valid,
      ins_ready => fork96_outs_0_ready,
      clk => clk,
      rst => rst,
      outs => extsi45_outs,
      outs_valid => extsi45_outs_valid,
      outs_ready => extsi45_outs_ready
    );

  extsi46 : entity work.extsi(arch) generic map(8, 11)
    port map(
      ins => fork96_outs_1,
      ins_valid => fork96_outs_1_valid,
      ins_ready => fork96_outs_1_ready,
      clk => clk,
      rst => rst,
      outs => extsi46_outs,
      outs_valid => extsi46_outs_valid,
      outs_ready => extsi46_outs_ready
    );

  extsi47 : entity work.extsi(arch) generic map(8, 11)
    port map(
      ins => fork96_outs_2,
      ins_valid => fork96_outs_2_valid,
      ins_ready => fork96_outs_2_ready,
      clk => clk,
      rst => rst,
      outs => extsi47_outs,
      outs_valid => extsi47_outs_valid,
      outs_ready => extsi47_outs_ready
    );

  cond_br261 : entity work.cond_br(arch) generic map(8)
    port map(
      condition => fork98_outs_6,
      condition_valid => fork98_outs_6_valid,
      condition_ready => fork98_outs_6_ready,
      data => cond_br258_falseOut,
      data_valid => cond_br258_falseOut_valid,
      data_ready => cond_br258_falseOut_ready,
      clk => clk,
      rst => rst,
      trueOut => cond_br261_trueOut,
      trueOut_valid => cond_br261_trueOut_valid,
      trueOut_ready => cond_br261_trueOut_ready,
      falseOut => cond_br261_falseOut,
      falseOut_valid => cond_br261_falseOut_valid,
      falseOut_ready => cond_br261_falseOut_ready
    );

  sink77 : entity work.sink(arch) generic map(8)
    port map(
      ins => cond_br261_falseOut,
      ins_valid => cond_br261_falseOut_valid,
      ins_ready => cond_br261_falseOut_ready,
      clk => clk,
      rst => rst
    );

  extsi48 : entity work.extsi(arch) generic map(8, 11)
    port map(
      ins => cond_br261_trueOut,
      ins_valid => cond_br261_trueOut_valid,
      ins_ready => cond_br261_trueOut_ready,
      clk => clk,
      rst => rst,
      outs => extsi48_outs,
      outs_valid => extsi48_outs_valid,
      outs_ready => extsi48_outs_ready
    );

  cond_br262 : entity work.cond_br(arch) generic map(32)
    port map(
      condition => fork98_outs_2,
      condition_valid => fork98_outs_2_valid,
      condition_ready => fork98_outs_2_ready,
      data => cond_br249_falseOut,
      data_valid => cond_br249_falseOut_valid,
      data_ready => cond_br249_falseOut_ready,
      clk => clk,
      rst => rst,
      trueOut => cond_br262_trueOut,
      trueOut_valid => cond_br262_trueOut_valid,
      trueOut_ready => cond_br262_trueOut_ready,
      falseOut => cond_br262_falseOut,
      falseOut_valid => cond_br262_falseOut_valid,
      falseOut_ready => cond_br262_falseOut_ready
    );

  sink78 : entity work.sink(arch) generic map(32)
    port map(
      ins => cond_br262_falseOut,
      ins_valid => cond_br262_falseOut_valid,
      ins_ready => cond_br262_falseOut_ready,
      clk => clk,
      rst => rst
    );

  cond_br263 : entity work.cond_br_dataless(arch)
    port map(
      condition => buffer272_outs,
      condition_valid => buffer272_outs_valid,
      condition_ready => buffer272_outs_ready,
      data_valid => cond_br257_falseOut_valid,
      data_ready => cond_br257_falseOut_ready,
      clk => clk,
      rst => rst,
      trueOut_valid => cond_br263_trueOut_valid,
      trueOut_ready => cond_br263_trueOut_ready,
      falseOut_valid => cond_br263_falseOut_valid,
      falseOut_ready => cond_br263_falseOut_ready
    );

  buffer272 : entity work.tfifo(arch) generic map(1, 1)
    port map(
      ins => fork98_outs_1,
      ins_valid => fork98_outs_1_valid,
      ins_ready => fork98_outs_1_ready,
      clk => clk,
      rst => rst,
      outs => buffer272_outs,
      outs_valid => buffer272_outs_valid,
      outs_ready => buffer272_outs_ready
    );

  sink79 : entity work.sink_dataless(arch)
    port map(
      ins_valid => cond_br263_falseOut_valid,
      ins_ready => cond_br263_falseOut_ready,
      clk => clk,
      rst => rst
    );

  extsi49 : entity work.extsi(arch) generic map(3, 4)
    port map(
      ins => cond_br8_falseOut,
      ins_valid => cond_br8_falseOut_valid,
      ins_ready => cond_br8_falseOut_ready,
      clk => clk,
      rst => rst,
      outs => extsi49_outs,
      outs_valid => extsi49_outs_valid,
      outs_ready => extsi49_outs_ready
    );

  source5 : entity work.source(arch)
    port map(
      clk => clk,
      rst => rst,
      outs_valid => source5_outs_valid,
      outs_ready => source5_outs_ready
    );

  constant29 : entity work.handshake_constant_5(arch) generic map(3)
    port map(
      ctrl_valid => source5_outs_valid,
      ctrl_ready => source5_outs_ready,
      clk => clk,
      rst => rst,
      outs => constant29_outs,
      outs_valid => constant29_outs_valid,
      outs_ready => constant29_outs_ready
    );

  extsi50 : entity work.extsi(arch) generic map(3, 4)
    port map(
      ins => constant29_outs,
      ins_valid => constant29_outs_valid,
      ins_ready => constant29_outs_ready,
      clk => clk,
      rst => rst,
      outs => extsi50_outs,
      outs_valid => extsi50_outs_valid,
      outs_ready => extsi50_outs_ready
    );

  source6 : entity work.source(arch)
    port map(
      clk => clk,
      rst => rst,
      outs_valid => source6_outs_valid,
      outs_ready => source6_outs_ready
    );

  constant30 : entity work.handshake_constant_2(arch) generic map(2)
    port map(
      ctrl_valid => source6_outs_valid,
      ctrl_ready => source6_outs_ready,
      clk => clk,
      rst => rst,
      outs => constant30_outs,
      outs_valid => constant30_outs_valid,
      outs_ready => constant30_outs_ready
    );

  extsi51 : entity work.extsi(arch) generic map(2, 4)
    port map(
      ins => constant30_outs,
      ins_valid => constant30_outs_valid,
      ins_ready => constant30_outs_ready,
      clk => clk,
      rst => rst,
      outs => extsi51_outs,
      outs_valid => extsi51_outs_valid,
      outs_ready => extsi51_outs_ready
    );

  addi6 : entity work.addi(arch) generic map(4)
    port map(
      lhs => extsi49_outs,
      lhs_valid => extsi49_outs_valid,
      lhs_ready => extsi49_outs_ready,
      rhs => extsi51_outs,
      rhs_valid => extsi51_outs_valid,
      rhs_ready => extsi51_outs_ready,
      clk => clk,
      rst => rst,
      result => addi6_result,
      result_valid => addi6_result_valid,
      result_ready => addi6_result_ready
    );

  buffer114 : entity work.oehb(arch) generic map(4)
    port map(
      ins => addi6_result,
      ins_valid => addi6_result_valid,
      ins_ready => addi6_result_ready,
      clk => clk,
      rst => rst,
      outs => buffer114_outs,
      outs_valid => buffer114_outs_valid,
      outs_ready => buffer114_outs_ready
    );

  fork97 : entity work.handshake_fork(arch) generic map(2, 4)
    port map(
      ins => buffer114_outs,
      ins_valid => buffer114_outs_valid,
      ins_ready => buffer114_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork97_outs_0,
      outs(1) => fork97_outs_1,
      outs_valid(0) => fork97_outs_0_valid,
      outs_valid(1) => fork97_outs_1_valid,
      outs_ready(0) => fork97_outs_0_ready,
      outs_ready(1) => fork97_outs_1_ready
    );

  trunci8 : entity work.trunci(arch) generic map(4, 3)
    port map(
      ins => fork97_outs_0,
      ins_valid => fork97_outs_0_valid,
      ins_ready => fork97_outs_0_ready,
      clk => clk,
      rst => rst,
      outs => trunci8_outs,
      outs_valid => trunci8_outs_valid,
      outs_ready => trunci8_outs_ready
    );

  cmpi2 : entity work.handshake_cmpi_2(arch) generic map(4)
    port map(
      lhs => fork97_outs_1,
      lhs_valid => fork97_outs_1_valid,
      lhs_ready => fork97_outs_1_ready,
      rhs => extsi50_outs,
      rhs_valid => extsi50_outs_valid,
      rhs_ready => extsi50_outs_ready,
      clk => clk,
      rst => rst,
      result => cmpi2_result,
      result_valid => cmpi2_result_valid,
      result_ready => cmpi2_result_ready
    );

  buffer115 : entity work.oehb(arch) generic map(1)
    port map(
      ins => cmpi2_result,
      ins_valid => cmpi2_result_valid,
      ins_ready => cmpi2_result_ready,
      clk => clk,
      rst => rst,
      outs => buffer115_outs,
      outs_valid => buffer115_outs_valid,
      outs_ready => buffer115_outs_ready
    );

  fork98 : entity work.handshake_fork(arch) generic map(8, 1)
    port map(
      ins => buffer115_outs,
      ins_valid => buffer115_outs_valid,
      ins_ready => buffer115_outs_ready,
      clk => clk,
      rst => rst,
      outs(0) => fork98_outs_0,
      outs(1) => fork98_outs_1,
      outs(2) => fork98_outs_2,
      outs(3) => fork98_outs_3,
      outs(4) => fork98_outs_4,
      outs(5) => fork98_outs_5,
      outs(6) => fork98_outs_6,
      outs(7) => fork98_outs_7,
      outs_valid(0) => fork98_outs_0_valid,
      outs_valid(1) => fork98_outs_1_valid,
      outs_valid(2) => fork98_outs_2_valid,
      outs_valid(3) => fork98_outs_3_valid,
      outs_valid(4) => fork98_outs_4_valid,
      outs_valid(5) => fork98_outs_5_valid,
      outs_valid(6) => fork98_outs_6_valid,
      outs_valid(7) => fork98_outs_7_valid,
      outs_ready(0) => fork98_outs_0_ready,
      outs_ready(1) => fork98_outs_1_ready,
      outs_ready(2) => fork98_outs_2_ready,
      outs_ready(3) => fork98_outs_3_ready,
      outs_ready(4) => fork98_outs_4_ready,
      outs_ready(5) => fork98_outs_5_ready,
      outs_ready(6) => fork98_outs_6_ready,
      outs_ready(7) => fork98_outs_7_ready
    );

  cond_br10 : entity work.cond_br(arch) generic map(3)
    port map(
      condition => fork98_outs_0,
      condition_valid => fork98_outs_0_valid,
      condition_ready => fork98_outs_0_ready,
      data => trunci8_outs,
      data_valid => trunci8_outs_valid,
      data_ready => trunci8_outs_ready,
      clk => clk,
      rst => rst,
      trueOut => cond_br10_trueOut,
      trueOut_valid => cond_br10_trueOut_valid,
      trueOut_ready => cond_br10_trueOut_ready,
      falseOut => cond_br10_falseOut,
      falseOut_valid => cond_br10_falseOut_valid,
      falseOut_ready => cond_br10_falseOut_ready
    );

  sink81 : entity work.sink(arch) generic map(3)
    port map(
      ins => cond_br10_falseOut,
      ins_valid => cond_br10_falseOut_valid,
      ins_ready => cond_br10_falseOut_ready,
      clk => clk,
      rst => rst
    );

  cond_br11 : entity work.cond_br_dataless(arch)
    port map(
      condition => buffer276_outs,
      condition_valid => buffer276_outs_valid,
      condition_ready => buffer276_outs_ready,
      data_valid => cond_br9_falseOut_valid,
      data_ready => cond_br9_falseOut_ready,
      clk => clk,
      rst => rst,
      trueOut_valid => cond_br11_trueOut_valid,
      trueOut_ready => cond_br11_trueOut_ready,
      falseOut_valid => cond_br11_falseOut_valid,
      falseOut_ready => cond_br11_falseOut_ready
    );

  buffer276 : entity work.tfifo(arch) generic map(1, 1)
    port map(
      ins => fork98_outs_5,
      ins_valid => fork98_outs_5_valid,
      ins_ready => fork98_outs_5_ready,
      clk => clk,
      rst => rst,
      outs => buffer276_outs,
      outs_valid => buffer276_outs_valid,
      outs_ready => buffer276_outs_ready
    );

  fork99 : entity work.fork_dataless(arch) generic map(2)
    port map(
      ins_valid => cond_br11_falseOut_valid,
      ins_ready => cond_br11_falseOut_ready,
      clk => clk,
      rst => rst,
      outs_valid(0) => fork99_outs_0_valid,
      outs_valid(1) => fork99_outs_1_valid,
      outs_ready(0) => fork99_outs_0_ready,
      outs_ready(1) => fork99_outs_1_ready
    );

end architecture;
