library IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;
use work.types.all;

entity specgenCore is
  generic (
    DATA_SIZE : integer
  );
  port (
    clk, rst : in std_logic;

    ins : in std_logic_vector(DATA_SIZE - 1 downto 0);
    ins_valid : in std_logic;
    ins_spec_tag : in std_logic;
    ins_ready : out std_logic;

    predict_ins : in std_logic_vector(DATA_SIZE - 1 downto 0);
    predict_ins_valid : in std_logic;
    predict_ins_ready : out std_logic;

    fifo_ins : in std_logic_vector(DATA_SIZE - 1 downto 0);
    fifo_ins_valid : in std_logic;
    fifo_ins_ready : out std_logic;

    outs : out std_logic_vector(DATA_SIZE - 1 downto 0);
    outs_spec_tag : out std_logic;

    fifo_outs : out std_logic_vector(DATA_SIZE - 1 downto 0);
    fifo_outs_valid : out std_logic;
    fifo_outs_ready : in std_logic;

    control_outs : out std_logic_vector(2 downto 0); -- 000:spec, 001:no cmp, 010:cmp correct, 011:resend, 100:kill, 101:correct-spec
    control_outs_valid : out std_logic;
    control_outs_ready : in std_logic
  );
end specgenCore;

architecture arch of specgenCore is

type State_type is (PASS, SPEC, NO_CMP, CMP_CORRECT, CMP_WRONG, KILL1, KILL2, KILL3, KILL_SPEC);
type Control_type is (CONTROL_SPEC, CONTROL_NO_CMP, CONTROL_CMP_CORRECT, CONTROL_RESEND, CONTROL_KILL, CONTROL_CORRECT_SPEC);
signal State : State_type;

signal DatapV : std_logic;
signal PredictpV : std_logic;
signal FifoNotEmpty : std_logic;
signal ControlnR : std_logic;
signal FifoNotFull : std_logic;

signal DataR : std_logic;
signal PredictR : std_logic;
signal FifoR : std_logic;
signal ControlV : std_logic;
signal FifoV : std_logic;

signal StateInternal : std_logic_vector(3 downto 0);
signal ControlInternal : Control_type;

begin
    DatapV <= ins_valid;
    PredictpV <= predict_ins_valid;
    FifoNotEmpty <= fifo_ins_valid;
    ControlnR <= control_outs_ready;
    FifoNotFull <= fifo_outs_ready;

    ins_ready <= DataR;
    predict_ins_ready <= PredictR;
    fifo_ins_ready <= FifoR;
    control_outs_valid <= ControlV;
    fifo_outs_valid <= FifoV;

process(ControlInternal)
    begin
        case ControlInternal is
            when CONTROL_SPEC =>
                control_outs <= "000";
            when CONTROL_NO_CMP =>
                control_outs <= "001";
            when CONTROL_CMP_CORRECT =>
                control_outs <= "010";
            when CONTROL_RESEND =>
                control_outs <= "011";
            when CONTROL_KILL =>
                control_outs <= "100";
            when CONTROL_CORRECT_SPEC =>
                control_outs <= "101";
        end case;
    end process;

process(State)
    begin
        case State is
            when PASS => -- 0
                StateInternal <= "0000";
            when SPEC => -- 1
                StateInternal <= "0001";
            when NO_CMP => -- 2
                StateInternal <= "0010";
            when CMP_CORRECT => -- 3
                StateInternal <= "0011";
            when CMP_WRONG => -- 4
                StateInternal <= "0100";
            when KILL1 => -- 5
                StateInternal <= "0101";
            when KILL2 => -- 6
                StateInternal <= "0110";
            when KILL3 => -- 7
                StateInternal <= "0111";
            when KILL_SPEC => -- 8
                StateInternal <= "1000";

        end case;

    end process;

state_proc : process (clk)
    begin
        if rising_edge(clk) then
            if rst = '1' then
                State <= PASS;
            else
                case State is
                    when PASS =>
                        if (DatapV = '0' and PredictpV = '1' and FifoNotFull = '1' and ControlnR = '0') then
                            State <= SPEC;
                        elsif (DatapV = '1' and FifoNotEmpty = '0' and ControlnR = '0') then
                            State <= NO_CMP;
                        elsif (DatapV = '1' and FifoNotEmpty = '1' and ins = fifo_ins and ControlnR = '0') then
                            State <= CMP_CORRECT;
                        elsif (DatapV = '1' and FifoNotEmpty = '1' and ins /= fifo_ins and ControlnR = '0') then
                            State <= CMP_WRONG;
                        elsif (DatapV = '1' and FifoNotEmpty = '1' and ins /= fifo_ins and ControlnR = '1') then
                            State <= KILL1;
                        end if;
                    when SPEC =>
                        if (ControlnR = '1') then
                            State <= PASS;
                        end if;
                    when NO_CMP =>
                        if (ControlnR = '1') then
                            State <= PASS;
                        end if;
                    when CMP_CORRECT =>
                        if (ControlnR = '1') then
                            State <= PASS;
                        end if;
                    when CMP_WRONG =>
                        if (ControlnR = '1') then
                            State <= KILL1;
                        end if;
                    when KILL1 =>
                        if (DatapV = '1' and ins_spec_tag = '0') then
                            if (FifoNotEmpty = '0') then
                                State <= PASS;
                            else
                                State <= KILL2;
                            end if;
                        elsif (FifoNotEmpty = '0') then
                            State <= KILL3;
                        end if;

                    when KILL2 =>
                        if (FifoNotEmpty = '0') then
                            State <= PASS;
                        end if;

                    when KILL3 =>
                        if ((DatapV = '0' or (DatapV = '1' and ins_spec_tag = '1')) and PredictpV = '1' and FifoNotFull = '1' and ControlnR = '0') then
                            State <= KILL_SPEC;
                        elsif (DatapV = '1' and ins_spec_tag = '0' and PredictpV = '1' and FifoNotFull = '1' and ControlnR = '0') then
                            State <= SPEC;
                        elsif (DatapV = '1' and ins_spec_tag = '0') then
                            State <= PASS;
                        end if;
                    when KILL_SPEC =>
                        if ((DatapV = '0' or (DatapV = '1' and ins_spec_tag = '1')) and ControlnR = '1') then
                            State <= KILL3;
                        elsif (DatapV = '1' and ins_spec_tag = '0' and ControlnR = '0') then
                            State <= SPEC;
                        elsif (DatapV = '1' and ins_spec_tag = '0' and ControlnR = '1') then
                            State <= PASS;
                        end if;
                end case;
            end if;
        end if;

    end process;

output_proc : process (State, ins, ins_spec_tag, fifo_ins, predict_ins, DatapV, PredictpV, FifoNotEmpty, ControlnR, FifoNotFull)
    begin

        outs <= ins;
        outs_spec_tag <= '0';
        fifo_outs <= predict_ins;
        ControlInternal <= CONTROL_SPEC;

        case State is
            when PASS =>
                DataR <= ControlnR;
                PredictR <= FifoNotFull and ControlnR;

                if (DatapV = '1' and FifoNotEmpty = '1' and ins = fifo_ins) then
                    FifoR <= '1';
                else
                    FifoR <= '0';
                end if;

                --FifoV <= not DatapV and PredictpV;
                FifoV <= '0';

                if (DatapV = '0' and PredictpV = '1' and FifoNotFull = '1') then
                    ControlV <= '1';
                    ControlInternal <= CONTROL_SPEC;
                    outs <= predict_ins;
                    outs_spec_tag <= '1';
                    FifoV <= '1';
                elsif (DatapV = '1' and FifoNotEmpty = '0') then
                    ControlV <= '1';
                    ControlInternal <= CONTROL_NO_CMP;
                    outs <= ins;
                    outs_spec_tag <= '0';
                elsif (DatapV = '1' and PredictpV = '1' and FifoNotEmpty = '1' and ins = fifo_ins) then
                    ControlV <= '1';
                    ControlInternal <= CONTROL_CORRECT_SPEC;
                    outs <= predict_ins;
                    outs_spec_tag <= '1';
                    FifoV <= '1';
                elsif (DatapV = '1' and PredictpV = '0' and FifoNotEmpty = '1' and ins = fifo_ins) then
                    ControlV <= '1';
                    ControlInternal <= CONTROL_CMP_CORRECT;
                elsif (DatapV = '1' and FifoNotEmpty = '1' and ins /= fifo_ins) then
                    ControlV <= '1';
                    ControlInternal <= CONTROL_RESEND;
                    outs <= ins;
                    outs_spec_tag <= '0';
                else
                    ControlV <= '0';
                end if;

            when SPEC =>
                DataR <= '0';
                PredictR <= ControlnR;
                FifoR <= '0';
                ControlV <= '1';
                FifoV <= '0';

                ControlInternal <= CONTROL_SPEC;

                outs <= predict_ins;
                outs_spec_tag <= '1';

            when NO_CMP =>
                DataR <= ControlnR;
                PredictR <= '0';
                FifoR <= '0';
                ControlV <= '1';
                FifoV <= '0';

                ControlInternal <= CONTROL_NO_CMP;

                outs <= ins;
                outs_spec_tag <= '0';

            when CMP_CORRECT =>
                DataR <= ControlnR;
                PredictR <= '0';
                FifoR <= '0';
                ControlV <= '1';
                FifoV <= '0';

                ControlInternal <= CONTROL_CMP_CORRECT;

            when CMP_WRONG =>
                DataR <= ControlnR;
                PredictR <= '0';
                FifoR <= '0';
                ControlV <= '1';
                FifoV <= '0';

                ControlInternal <= CONTROL_RESEND;

                outs <= ins;
                outs_spec_tag <= '0';

            when KILL1 =>
                DataR <= DatapV and ins_spec_tag;
                FifoR <= ControlnR;
                PredictR<= '0';
                ControlV <= FifoNotEmpty;
                FifoV <= '0';

                ControlInternal <= CONTROL_KILL;

            when KILL2 =>
                DataR <= '0';
                FifoR <= ControlnR;
                PredictR<= '0';
                ControlV <= FifoNotEmpty;
                FifoV <= '0';

                ControlInternal <= CONTROL_KILL;

            when KILL3 =>
                DataR <= DatapV and ins_spec_tag;
                PredictR <= ControlnR;
                FifoR <= '0';
                ControlV <= PredictpV and FifoNotFull;
                FifoV <= PredictpV;

                ControlInternal <= CONTROL_SPEC;

                outs <= predict_ins;
                outs_spec_tag <= '1';

            when KILL_SPEC =>
                DataR <= DatapV and ins_spec_tag;
                PredictR <= ControlnR;
                FifoR <= '0';
                ControlV <= '1';
                FifoV <= '0';

                ControlInternal <= CONTROL_SPEC;

                outs <= predict_ins;
                outs_spec_tag <= '1';

        end case;

    end process;

end architecture;


library IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;
use work.types.all;
entity decodeSave is
  port (
    control_in : in std_logic_vector(2 downto 0);
    control_in_valid : in std_logic;
    control_in_ready : out std_logic;

    control_out : out std_logic_vector(0 downto 0); -- 0:resend, 1:drop
    control_out_valid : out std_logic;
    control_out_ready : in std_logic
  );
end decodeSave;

architecture arch of decodeSave is

begin
    process (control_in, control_in_valid, control_out_ready)
    begin
        if (control_in = "001" or control_in = "010" or control_in = "011" or control_in = "101") then
            control_in_ready <= control_out_ready;
        else
            control_in_ready <= '1';
        end if;

        control_out_valid <= '0';
        control_out(0) <= '0';

        if (control_in_valid = '1') then
            if control_in = "001" then -- no cmp
                control_out_valid <= '1';
                control_out(0) <= '1';
            elsif control_in = "010" then -- cmp correct
                control_out_valid <= '1';
                control_out(0) <= '1';
            elsif control_in = "101" then -- correct-spec
                control_out_valid <= '1';
                control_out(0) <= '1';
            elsif control_in = "011" then --cmp wrong
                control_out_valid <= '1';
                control_out(0) <= '0';
            end if;
        end if;

    end process;
end architecture;


library IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;
use work.types.all;
entity decodeCommit is
  port (
    control_in : in std_logic_vector(2 downto 0);
    control_in_valid : in std_logic;
    control_in_ready : out std_logic;

    control_out : out std_logic_vector(0 downto 0); -- 0:pass, 1:discard
    control_out_valid : out std_logic;
    control_out_ready : in std_logic
  );
end decodeCommit;

architecture arch of decodeCommit is

begin
    process (control_in, control_in_valid, control_out_ready)
    begin
        if (control_in = "010" or control_in = "100" or control_in = "101") then
            control_in_ready <= control_out_ready;
        else
            control_in_ready <= '1';
        end if;

        control_out_valid <= '0';
        control_out(0) <= '0';

        if (control_in_valid = '1') then
            if control_in = "010" then -- cmp correct
                control_out_valid <= '1';
                control_out(0) <= '0';
            elsif control_in = "101" then -- correct-spec
                control_out_valid <= '1';
                control_out(0) <= '0';
            elsif control_in = "100" then -- cmp wrong
                control_out_valid <= '1';
                control_out(0) <= '1';
            end if;
        end if;

    end process;
end architecture;



library IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;
use work.types.all;
entity decodeBranch is
  port (
    control_in : in std_logic_vector(2 downto 0);
    control_in_valid : in std_logic;
    control_in_ready : out std_logic;

    control_out : out std_logic_vector(0 downto 0); -- 1:pass, 0:discard
    control_out_valid : out std_logic;
    control_out_ready : in std_logic
  );
end decodeBranch;

architecture arch of decodeBranch is

begin
    process (control_in, control_in_valid, control_out_ready)
    begin
        if (control_in = "010" or control_in = "100" or control_in = "101") then
            control_in_ready <= control_out_ready;
        else
            control_in_ready <= '1';
        end if;

        control_out_valid <= '0';
        control_out(0) <= '0';

        if (control_in_valid = '1') then
            if control_in = "010" then -- cmp correct
                control_out_valid <= '1';
                control_out(0) <= '0';
            elsif control_in = "101" then -- correct-spec
                control_out_valid <= '1';
                control_out(0) <= '0';
            elsif control_in = "100" then --cmp wrong
                control_out_valid <= '1';
                control_out(0) <= '1';
            end if;
        end if;

    end process;
end architecture;



library IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;
use work.types.all;
entity decodeSC is
  port (
    control_in : in std_logic_vector(2 downto 0);
    control_in_valid : in std_logic;
    control_in_ready : out std_logic;

    control_out0 : out std_logic_vector(2 downto 0); -- 000:pass, 001:kill, 010:resend, 011:kill-pass, 100:no_cmp
    control_out0_valid : out std_logic;
    control_out0_ready : in std_logic;

    control_out1 : out std_logic_vector(2 downto 0); -- 000:pass, 001:kill, 010:resend, 011:kill-pass, 100:no_cmp
    control_out1_valid : out std_logic;
    control_out1_ready : in std_logic
  );
end decodeSC;

architecture arch of decodeSC is

begin
    process (control_in, control_in_valid, control_out0_ready, control_out1_ready)
    begin
        if (control_in = "000" or control_in = "001" or control_in = "010" or control_in = "011" or control_in = "101") then
            control_in_ready <= control_out0_ready;
        else
            control_in_ready <= control_out1_ready;
        end if;

        control_out0_valid <= '0';
        control_out1_valid <= '0';
        control_out0 <= "000";
        control_out1 <= "000";

        if (control_in_valid = '1') then
            if control_in = "000" then -- spec
                control_out0_valid <= '1';
                control_out0 <= "000";
            elsif control_in = "001" then -- no cmp
                control_out0_valid <= '1';
                control_out0 <= "100";
            elsif control_in = "010" then -- cmp correct
                control_out0_valid <= '1';
                control_out0 <= "001";
            elsif control_in = "101" then -- correct-spec
                control_out0_valid <= '1';
                control_out0 <= "011";
            elsif control_in = "011" then -- cmp wrong resend
                control_out0_valid <= '1';
                control_out0 <= "010";
            elsif control_in = "100" then -- cmp wrong kill
                control_out1_valid <= '1';
                control_out1 <= "001";
            end if;
        end if;

    end process;
end architecture;

library IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;
use work.types.all;
entity decodeOutput is
  port (
    control_in : in std_logic_vector(2 downto 0);
    control_in_valid : in std_logic;
    control_in_ready : out std_logic;

    out_valid : out std_logic;
    out_ready : in std_logic
  );
end decodeOutput;

architecture arch of decodeOutput is

begin
    process (control_in, control_in_valid, out_ready)
    begin
        if (control_in = "000" or control_in = "001" or control_in = "011" or control_in = "101") then
            control_in_ready <= out_ready;
        else
            control_in_ready <= '1';
        end if;

        out_valid <= '0';

        if (control_in_valid = '1') then
            if control_in = "000" then -- spec
                out_valid <= '1';
            elsif control_in = "101" then -- correct-spec
                out_valid <= '1';
            elsif control_in = "001" then -- no cmp
                out_valid <= '1';
            elsif control_in = "011" then -- cmp wrong resend
                out_valid <= '1';
            end if;
        end if;

    end process;
end architecture;


library IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;
use work.types.all;
entity predictor is
  generic (
    DATA_SIZE : integer -- use normal data size, eg- 32
  );
  port (
    clk, rst     : in  std_logic;

    enable_valid : in std_logic;
    enable_ready : out std_logic;

    data_in      : in std_logic_vector(DATA_SIZE - 1 downto 0);
    data_in_valid : in std_logic;
    data_in_ready : out std_logic;

    data_out     : out std_logic_vector(DATA_SIZE - 1 downto 0);
    data_out_valid : out std_logic;
    data_out_ready : in std_logic
  );
end predictor;

architecture arch of predictor is
    signal zeros : std_logic_vector(DATA_SIZE-2 downto 0);
    signal data_reg: std_logic_vector(DATA_SIZE-1 downto 0);

begin

    zeros <= (others => '0');

    --predicted value is 1 by default and updated to the latest real value
    process(clk, rst) is
          begin
           if (rst = '1') then

            data_reg <= zeros & '1';

            elsif (rising_edge(clk)) then
                if (data_in_valid = '1') then
                    data_reg <= data_in;
                end if;
            end if;
    end process;

    enable_ready <= data_out_ready;
    data_in_ready <= data_out_ready;

    -- Predictor output valid if enabled
    data_out <= data_reg; -- zeros & '1';
    data_out_valid <= enable_valid;
end arch;

library IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;
use work.types.all;

entity predFifo is
  generic (
    DATA_SIZE : integer;
    FIFO_DEPTH : integer
  );
  port (
    clk, rst : in std_logic;

    data_in : in std_logic_vector(DATA_SIZE - 1 downto 0);
    data_in_valid : in std_logic;
    data_in_ready : out std_logic;

    data_out : out std_logic_vector(DATA_SIZE - 1 downto 0);
    data_out_valid : out std_logic;
    data_out_ready : in std_logic
  );
end predFifo;

architecture arch of predFifo is

    signal HeadEn   : std_logic := '0';
    signal TailEn  : std_logic := '0';

    signal Tail : natural range 0 to FIFO_DEPTH - 1;
    signal Head : natural range 0 to FIFO_DEPTH - 1;

    signal Empty    : std_logic;
    signal Full : std_logic;

    type FIFO_Memory is array (0 to FIFO_DEPTH - 1) of STD_LOGIC_VECTOR (DATA_SIZE-1 downto 0);
    signal Memory : FIFO_Memory;


begin
    data_out_valid <= not Empty;
    data_in_ready <= not Full;

    TailEn <= not Full and data_in_valid;
    HeadEn <= not Empty and data_out_ready;
    data_out <= Memory(Head);

----------------------------------------------------------------

-- Sequential Process

----------------------------------------------------------------

-------------------------------------------
-- process for writing data
fifo_proc : process (clk)

     begin
        if rising_edge(clk) then
          if rst = '1' then

          else

            if (TailEn = '1' ) then
                -- Write Data to Memory
                Memory(Tail) <= data_in;

            end if;

          end if;
        end if;
    end process;



-------------------------------------------
-- process for updating tail
TailUpdate_proc : process (clk)

      begin
        if rising_edge(clk) then

            if rst = '1' then
               Tail <= 0;
            else

                if (TailEn = '1') then

                    Tail  <= (Tail + 1) mod FIFO_DEPTH;

                end if;

            end if;
        end if;
    end process;

-------------------------------------------
-- process for updating head
HeadUpdate_proc : process (clk)

  begin
  if rising_edge(clk) then

    if rst = '1' then
       Head <= 0;
    else

        if (HeadEn = '1') then

            Head  <= (Head + 1) mod FIFO_DEPTH;

        end if;

    end if;
  end if;
end process;

-------------------------------------------
-- process for updating full
FullUpdate_proc : process (clk)

  begin
  if rising_edge(clk) then

    if rst = '1' then
       Full <= '0';
    else

        -- if only filling but not emptying
        if (TailEn = '1') and (HeadEn = '0') then

            -- if new tail index will reach head index
            if ((Tail +1) mod FIFO_DEPTH = Head) then

                Full  <= '1';

            end if;
        -- if only emptying but not filling
        elsif (TailEn = '0') and (HeadEn = '1') then
                Full <= '0';
        -- otherwise, nothing is happening or simultaneous read and write

        end if;

    end if;
  end if;
end process;

 -------------------------------------------
-- process for updating empty
EmptyUpdate_proc : process (clk)

  begin
  if rising_edge(clk) then

    if rst = '1' then
       Empty <= '1';
    else
        -- if only emptying but not filling
        if (TailEn = '0') and (HeadEn = '1') then

            -- if new head index will reach tail index
            if ((Head +1) mod FIFO_DEPTH = Tail) then

                Empty  <= '1';

            end if;
        -- if only filling but not emptying
        elsif (TailEn = '1') and (HeadEn = '0') then
                Empty <= '0';
       -- otherwise, nothing is happening or simultaneous read and write

        end if;

    end if;
  end if;
end process;

end architecture;

library ieee;
use ieee.std_logic_1164.all;
use work.types.all;
entity speculator is
  generic (
    DATA_TYPE : integer; -- use normal data size, eg- 32
    FIFO_DEPTH    : integer -- extra parameter for FIFO
  );
  port (
    clk, rst : in  std_logic;
    -- inputs
    ins: in std_logic_vector(DATA_TYPE - 1 downto 0);
    ins_valid: in std_logic;
    ins_spec_tag: in std_logic;
    ins_ready: out std_logic;
    -- enable is dataless (control token)
    enable_valid: in std_logic;
    enable_spec_tag: in std_logic;
    enable_ready: out std_logic;
    -- outputs
    outs: out std_logic_vector(DATA_TYPE - 1 downto 0);
    outs_valid: out std_logic;
    outs_spec_tag: out std_logic;
    outs_ready: in std_logic;
    -- control signals
    ctrl_save: out std_logic_vector(0 downto 0);
    ctrl_save_valid: out std_logic;
    ctrl_save_spec_tag: out std_logic;
    ctrl_save_ready: in std_logic;
    ctrl_commit: out std_logic_vector(0 downto 0);
    ctrl_commit_valid: out std_logic;
    ctrl_commit_spec_tag: out std_logic;
    ctrl_commit_ready: in std_logic;
    ctrl_sc_save: out std_logic_vector(2 downto 0);
    ctrl_sc_save_valid: out std_logic;
    ctrl_sc_save_spec_tag: out std_logic;
    ctrl_sc_save_ready: in std_logic;
    ctrl_sc_commit: out std_logic_vector(2 downto 0);
    ctrl_sc_commit_valid: out std_logic;
    ctrl_sc_commit_spec_tag: out std_logic;
    ctrl_sc_commit_ready: in std_logic;
    ctrl_sc_branch: out std_logic_vector(0 downto 0);
    ctrl_sc_branch_valid: out std_logic;
    ctrl_sc_branch_spec_tag: out std_logic;
    ctrl_sc_branch_ready: in std_logic
  );
end speculator;

architecture arch of speculator is
signal fork_data_outs : data_array (1 downto 0)(DATA_TYPE - 1 downto 0);
signal fork_data_outs_valid : std_logic_vector(1 downto 0);
signal fork_data_outs_spec_tag : std_logic_vector(1 downto 0);
signal fork_data_outs_ready : std_logic_vector(1 downto 0);

signal predictor_data_out : std_logic_vector(DATA_TYPE - 1 downto 0);
signal predictor_data_out_valid : std_logic;
signal predictor_data_out_ready : std_logic;

signal specgenCore_fifo_outs : std_logic_vector(DATA_TYPE - 1 downto 0);
signal specgenCore_fifo_outs_valid : std_logic;
signal specgenCore_fifo_outs_ready : std_logic;

signal specgenCore_control_outs : std_logic_vector(2 downto 0);
signal specgenCore_control_outs_valid : std_logic;
signal specgenCore_control_outs_ready : std_logic;

signal predFifo_data_out : std_logic_vector(DATA_TYPE - 1 downto 0);
signal predFifo_data_out_valid : std_logic;
signal predFifo_data_out_ready : std_logic;

signal fork_control_outs : data_array (4 downto 0)(2 downto 0);
signal fork_control_outs_valid : std_logic_vector(4 downto 0);
signal fork_control_outs_ready : std_logic_vector(4 downto 0);
begin

ctrl_save_spec_tag <= '0';
ctrl_commit_spec_tag <= '0';
ctrl_sc_save_spec_tag <= '0';
ctrl_sc_commit_spec_tag <= '0';
ctrl_sc_branch_spec_tag <= '0';

data_fork: entity work.handshake_fork_with_tag(arch)
  generic map(
    SIZE => 2,
    DATA_TYPE => DATA_TYPE
  )
  port map(
    clk => clk,
    rst => rst,
    ins => ins,
    ins_valid => ins_valid,
    ins_spec_tag => ins_spec_tag,
    ins_ready => ins_ready,
    outs => fork_data_outs,
    outs_valid => fork_data_outs_valid,
    outs_spec_tag => fork_data_outs_spec_tag,
    outs_ready => fork_data_outs_ready
  );

spengenCore0: entity work.specgenCore(arch)
  generic map(
    DATA_SIZE => DATA_TYPE
  )
  port map (
    clk => clk,
    rst => rst,

    ins => fork_data_outs(0),
    ins_valid => fork_data_outs_valid(0),
    ins_spec_tag => fork_data_outs_spec_tag(0),
    ins_ready => fork_data_outs_ready(0),

    predict_ins => predictor_data_out,
    predict_ins_valid => predictor_data_out_valid,
    predict_ins_ready => predictor_data_out_ready,

    fifo_ins => predFifo_data_out,
    fifo_ins_valid => predFifo_data_out_valid,
    fifo_ins_ready => predFifo_data_out_ready,

    outs => outs,
    outs_spec_tag => outs_spec_tag,

    fifo_outs => specgenCore_fifo_outs,
    fifo_outs_valid => specgenCore_fifo_outs_valid,
    fifo_outs_ready => specgenCore_fifo_outs_ready,

    control_outs => specgenCore_control_outs,
    control_outs_valid => specgenCore_control_outs_valid,
    control_outs_ready => specgenCore_control_outs_ready
  );

predictor0: entity work.predictor(arch)
  generic map(
    DATA_SIZE => DATA_TYPE
  )
  port map (
    clk => clk,
    rst => rst,

    enable_valid => enable_valid,
    enable_ready => enable_ready,

    data_in => fork_data_outs(1),
    data_in_valid => fork_data_outs_valid(1),
    data_in_ready => fork_data_outs_ready(1),

    data_out => predictor_data_out,
    data_out_valid => predictor_data_out_valid,
    data_out_ready => predictor_data_out_ready
  );

predFifo0: entity work.predFifo(arch)
  generic map(
    DATA_SIZE => DATA_TYPE,
    FIFO_DEPTH => FIFO_DEPTH
  )
  port map (
    clk => clk,
    rst => rst,

    data_in => specgenCore_fifo_outs,
    data_in_valid => specgenCore_fifo_outs_valid,
    data_in_ready => specgenCore_fifo_outs_ready,

    data_out => predFifo_data_out,
    data_out_valid => predFifo_data_out_valid,
    data_out_ready => predFifo_data_out_ready
  );

fork0: entity work.handshake_fork(arch)
  generic map(
    SIZE => 5,
    DATA_TYPE => 3
  )
  port map (
    clk => clk,
    rst => rst,
    ins => specgenCore_control_outs,
    ins_valid => specgenCore_control_outs_valid,
    ins_ready => specgenCore_control_outs_ready,
    outs => fork_control_outs,
    outs_valid => fork_control_outs_valid,
    outs_ready => fork_control_outs_ready
  );

decodeSave0: entity work.decodeSave(arch)
  port map (
    control_in => fork_control_outs(3),
    control_in_valid => fork_control_outs_valid(3),
    control_in_ready => fork_control_outs_ready(3),
    control_out => ctrl_save,
    control_out_valid => ctrl_save_valid,
    control_out_ready => ctrl_save_ready
  );

decodeCommit0: entity work.decodeCommit(arch)
  port map (
    control_in => fork_control_outs(2),
    control_in_valid => fork_control_outs_valid(2),
    control_in_ready => fork_control_outs_ready(2),
    control_out => ctrl_commit,
    control_out_valid => ctrl_commit_valid,
    control_out_ready => ctrl_commit_ready
);

decodeSC0: entity work.decodeSC(arch)
  port map (
    control_in => fork_control_outs(1),
    control_in_valid => fork_control_outs_valid(1),
    control_in_ready => fork_control_outs_ready(1),
    control_out0 => ctrl_sc_save,
    control_out0_valid => ctrl_sc_save_valid,
    control_out0_ready => ctrl_sc_save_ready,
    control_out1 => ctrl_sc_commit,
    control_out1_valid => ctrl_sc_commit_valid,
    control_out1_ready => ctrl_sc_commit_ready
  );

decodeOutput0: entity work.decodeOutput(arch)
  port map (
    control_in => fork_control_outs(4),
    control_in_valid => fork_control_outs_valid(4),
    control_in_ready => fork_control_outs_ready(4),
    out_valid => outs_valid,
    out_ready => outs_ready
  );

decodeBranch0: entity work.decodeBranch(arch)
  port map (
    control_in => fork_control_outs(0),
    control_in_valid => fork_control_outs_valid(0),
    control_in_ready => fork_control_outs_ready(0),
    control_out => ctrl_sc_branch,
    control_out_valid => ctrl_sc_branch_valid,
    control_out_ready => ctrl_sc_branch_ready
  );
end arch;
