library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity cond_br_dataless is
  port (
    clk, rst : in std_logic;
    -- data input channel
    data_valid : in  std_logic;
    data_ready : out std_logic;
    -- condition input channel
    condition       : in  std_logic_vector(0 downto 0);
    condition_valid : in  std_logic;
    condition_ready : out std_logic;
    -- true output channel
    trueOut_valid : out std_logic;
    trueOut_ready : in  std_logic;
    -- false output channel
    falseOut_valid : out std_logic;
    falseOut_ready : in  std_logic
  );
end entity;

architecture arch of cond_br_dataless is
  signal joinValid, brReady : std_logic;
begin

  j : entity work.join(arch) generic map(2)
    port map(
    ins_valid(0) => data_valid,
    ins_valid(1) => condition_valid,
    outs_ready => brReady,
    outs_valid => joinValid,
    ins_ready(0) => data_ready, 
    ins_ready(1) => condition_ready);

  cond_brp : entity work.branch_simple(arch)
    port map(
      condition => condition(0),
      valid => joinValid,
      trueOut_ready => trueOut_ready,
      falseOut_ready => falseOut_ready,
      trueOut_valid => trueOut_valid,
      falseOut_valid => falseOut_valid,
      ins_ready => brReady);
end architecture;
