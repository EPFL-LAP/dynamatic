library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity ENTITY_NAME is
  generic (
    BITWIDTH : integer
  );
  port (
    -- inputs
    clk        : in std_logic;
    rst        : in std_logic;
    ctrl       : in std_logic_vector(0 downto 0);
    ctrl_valid : in std_logic;
    outs_ready : in std_logic;
    -- outputs
    ctrl_ready : out std_logic;
    outs       : out std_logic_vector(BITWIDTH - 1 downto 0);
    outs_valid : out std_logic);
end entity;

architecture arch of ENTITY_NAME is
begin
  outs       <= "VALUE";
  outs_valid <= ctrl_valid;
  ctrl_ready <= outs_ready;
end architecture;
