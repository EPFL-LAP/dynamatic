module __xls_float_ips__addf32_0_next(
  input wire clk,
  input wire rst,
  input wire [31:0] xls_float_ips__rhs,
  input wire xls_float_ips__rhs_vld,
  input wire [31:0] xls_float_ips__lhs,
  input wire xls_float_ips__lhs_vld,
  input wire xls_float_ips__result_rdy,
  output wire [31:0] xls_float_ips__result,
  output wire xls_float_ips__result_vld,
  output wire xls_float_ips__rhs_rdy,
  output wire xls_float_ips__lhs_rdy
);
  function automatic [3:0] priority_sel_4b_2way (input reg [1:0] sel, input reg [3:0] case0, input reg [3:0] case1, input reg [3:0] default_value);
    begin
      casez (sel)
        2'b?1: begin
          priority_sel_4b_2way = case0;
        end
        2'b10: begin
          priority_sel_4b_2way = case1;
        end
        2'b00: begin
          priority_sel_4b_2way = default_value;
        end
        default: begin
          // Propagate X
          priority_sel_4b_2way = 4'dx;
        end
      endcase
    end
  endfunction
  function automatic [1:0] priority_sel_2b_2way (input reg [1:0] sel, input reg [1:0] case0, input reg [1:0] case1, input reg [1:0] default_value);
    begin
      casez (sel)
        2'b?1: begin
          priority_sel_2b_2way = case0;
        end
        2'b10: begin
          priority_sel_2b_2way = case1;
        end
        2'b00: begin
          priority_sel_2b_2way = default_value;
        end
        default: begin
          // Propagate X
          priority_sel_2b_2way = 2'dx;
        end
      endcase
    end
  endfunction
  function automatic priority_sel_1b_4way (input reg [3:0] sel, input reg case0, input reg case1, input reg case2, input reg case3, input reg default_value);
    begin
      casez (sel)
        4'b???1: begin
          priority_sel_1b_4way = case0;
        end
        4'b??10: begin
          priority_sel_1b_4way = case1;
        end
        4'b?100: begin
          priority_sel_1b_4way = case2;
        end
        4'b1000: begin
          priority_sel_1b_4way = case3;
        end
        4'b0000: begin
          priority_sel_1b_4way = default_value;
        end
        default: begin
          // Propagate X
          priority_sel_1b_4way = 1'dx;
        end
      endcase
    end
  endfunction
  function automatic priority_sel_1b_3way (input reg [2:0] sel, input reg case0, input reg case1, input reg case2, input reg default_value);
    begin
      casez (sel)
        3'b??1: begin
          priority_sel_1b_3way = case0;
        end
        3'b?10: begin
          priority_sel_1b_3way = case1;
        end
        3'b100: begin
          priority_sel_1b_3way = case2;
        end
        3'b000: begin
          priority_sel_1b_3way = default_value;
        end
        default: begin
          // Propagate X
          priority_sel_1b_3way = 1'dx;
        end
      endcase
    end
  endfunction
  function automatic [2:0] priority_sel_3b_2way (input reg [1:0] sel, input reg [2:0] case0, input reg [2:0] case1, input reg [2:0] default_value);
    begin
      casez (sel)
        2'b?1: begin
          priority_sel_3b_2way = case0;
        end
        2'b10: begin
          priority_sel_3b_2way = case1;
        end
        2'b00: begin
          priority_sel_3b_2way = default_value;
        end
        default: begin
          // Propagate X
          priority_sel_3b_2way = 3'dx;
        end
      endcase
    end
  endfunction
  function automatic [1:0] priority_sel_2b_4way (input reg [3:0] sel, input reg [1:0] case0, input reg [1:0] case1, input reg [1:0] case2, input reg [1:0] case3, input reg [1:0] default_value);
    begin
      casez (sel)
        4'b???1: begin
          priority_sel_2b_4way = case0;
        end
        4'b??10: begin
          priority_sel_2b_4way = case1;
        end
        4'b?100: begin
          priority_sel_2b_4way = case2;
        end
        4'b1000: begin
          priority_sel_2b_4way = case3;
        end
        4'b0000: begin
          priority_sel_2b_4way = default_value;
        end
        default: begin
          // Propagate X
          priority_sel_2b_4way = 2'dx;
        end
      endcase
    end
  endfunction
  function automatic priority_sel_1b_2way (input reg [1:0] sel, input reg case0, input reg case1, input reg default_value);
    begin
      casez (sel)
        2'b?1: begin
          priority_sel_1b_2way = case0;
        end
        2'b10: begin
          priority_sel_1b_2way = case1;
        end
        2'b00: begin
          priority_sel_1b_2way = default_value;
        end
        default: begin
          // Propagate X
          priority_sel_1b_2way = 1'dx;
        end
      endcase
    end
  endfunction
  wire [31:0] __xls_float_ips__result_reg_init = {1'h0, 8'h00, 23'h00_0000};
  reg [7:0] p0_b_bexp__5;
  reg [7:0] p0_a_bexp__1;
  reg p0_bit_slice_92360;
  reg [22:0] p0_tuple_index_92361;
  reg [22:0] p0_tuple_index_92362;
  reg [7:0] p0_bit_slice_92363;
  reg p0_tuple_index_92364;
  reg p0_tuple_index_92365;
  reg [7:0] p1_a_bexp;
  reg p1_b_sign;
  reg p1_xor_92419;
  reg [24:0] p1_wide_x_squeezed;
  reg [24:0] p1_bit_slice_92421;
  reg [27:0] p1_shrl_92422;
  reg p1_sticky;
  reg p1_is_operand_inf;
  reg p1_and_92452;
  reg p1_is_result_nan;
  reg p1_not_92454;
  reg [7:0] p2_a_bexp;
  reg [27:0] p2_abs_fraction;
  reg p2_not_92500;
  reg p2_is_operand_inf;
  reg p2_is_result_nan;
  reg p2_result_sign;
  reg p2_not_92454;
  reg [7:0] p3_a_bexp;
  reg [27:0] p3_abs_fraction;
  reg p3_carry_bit;
  reg p3_and_92641;
  reg p3_and_92643;
  reg p3_nor_92649;
  reg p3_nor_92676;
  reg p3_leading_zeroes__4_to_5;
  reg [2:0] p3_priority_sel_92678;
  reg [1:0] p3_priority_sel_92679;
  reg [2:0] p3_priority_sel_92680;
  reg p3_or_92681;
  reg p3_not_92500;
  reg p3_is_operand_inf;
  reg p3_is_result_nan;
  reg p3_result_sign__2;
  reg [7:0] p4_a_bexp;
  reg p4_leading_zeroes__4_to_5;
  reg [3:0] p4_leading_zeroes__0_to_4;
  reg [2:0] p4_normal_chunk;
  reg [1:0] p4_half_way_chunk;
  reg [23:0] p4_bit_slice_92735;
  reg p4_not_92500;
  reg p4_is_operand_inf;
  reg p4_is_result_nan;
  reg p4_result_sign__2;
  reg p5_leading_zeroes__4_to_5;
  reg [3:0] p5_leading_zeroes__0_to_4;
  reg [9:0] p5_concat_92775;
  reg p5_not_92500;
  reg p5_is_operand_inf;
  reg p5_is_result_nan;
  reg [22:0] p5_result_fraction;
  reg p5_result_sign__2;
  reg [8:0] p6_wide_exponent__2;
  reg p6_is_operand_inf;
  reg p6_is_result_nan;
  reg [22:0] p6_result_fraction;
  reg p6_result_sign__2;
  reg p7_is_result_nan;
  reg [22:0] p7_result_fraction__3;
  reg p7_result_sign__2;
  reg [7:0] p7_result_exponent__2;
  reg p0_valid;
  reg p1_valid;
  reg p2_valid;
  reg p3_valid;
  reg p4_valid;
  reg p5_valid;
  reg p6_valid;
  reg p7_valid;
  reg [31:0] __xls_float_ips__result_reg;
  reg __xls_float_ips__result_valid_reg;
  wire xls_float_ips__result_valid_inv;
  wire xls_float_ips__result_valid_load_en;
  wire xls_float_ips__result_load_en;
  wire p8_stage_done;
  wire p8_not_valid;
  wire p7_enable;
  wire p7_data_enable;
  wire p7_not_valid;
  wire p6_enable;
  wire p6_data_enable;
  wire p6_not_valid;
  wire p5_enable;
  wire p5_data_enable;
  wire p5_not_valid;
  wire p4_enable;
  wire p4_data_enable;
  wire p4_not_valid;
  wire [2:0] fraction_shift__3;
  wire p3_enable;
  wire [9:0] add_92802;
  wire [24:0] concat_92763;
  wire carry_bit;
  wire [24:0] addend_x__1_squeezed;
  wire [7:0] a_bexp;
  wire [7:0] incremented_sum__1;
  wire [7:0] MAX_EXPONENT;
  wire [22:0] a_fraction;
  wire [7:0] b_bexp;
  wire [7:0] MAX_EXPONENT__1;
  wire [22:0] b_fraction;
  wire p3_data_enable;
  wire p3_not_valid;
  wire [9:0] wide_exponent;
  wire do_round_up;
  wire [24:0] add_92766;
  wire [3:0] leading_zeroes__0_to_4;
  wire nor_92548;
  wire nor_92549;
  wire nor_92551;
  wire nor_92552;
  wire nor_92557;
  wire nor_92558;
  wire nor_92563;
  wire nor_92566;
  wire nor_92567;
  wire nor_92568;
  wire nor_92574;
  wire [7:0] a_bexpbs_difference__1;
  wire eq_92432;
  wire eq_92433;
  wire eq_92434;
  wire eq_92435;
  wire p2_enable;
  wire and_reduce_92829;
  wire [9:0] wide_exponent__1;
  wire [24:0] rounded_fraction_squeezed_portion_3_width_25;
  wire [4:0] leading_zeroes;
  wire nor_92575;
  wire and_92576;
  wire and_92578;
  wire nor_92583;
  wire and_92584;
  wire nor_92587;
  wire and_92591;
  wire nor_92592;
  wire and_92596;
  wire nor_92598;
  wire [25:0] add_92484;
  wire [23:0] fraction_x;
  wire a_sign;
  wire b_sign;
  wire p2_data_enable;
  wire p2_not_valid;
  wire [7:0] b_bexp__5;
  wire rounding_carry;
  wire [2:0] fraction_shift__2;
  wire [2:0] fraction_shift__4;
  wire [28:0] cancel_fraction;
  wire and_92605;
  wire and_92623;
  wire [23:0] fraction_x__1;
  wire [2:0] addend_x__1_squeezed_const_lsb_bits__1;
  wire [23:0] fraction_y;
  wire [23:0] sign_ext_92404;
  wire [27:0] add_92423;
  wire p1_enable;
  wire [7:0] a_bexp__1;
  wire [27:0] rounded_fraction;
  wire [2:0] fraction_shift__1;
  wire [26:0] cancel_fraction__1;
  wire [26:0] carry_fraction__1;
  wire and_92641;
  wire and_92643;
  wire nor_92649;
  wire and_92650;
  wire [1:0] priority_sel_92657;
  wire [27:0] concat_92489;
  wire fraction_is_zero;
  wire [27:0] wide_x;
  wire [23:0] fraction_y__1;
  wire [2:0] addend_x__1_squeezed_const_lsb_bits;
  wire has_pos_inf;
  wire has_neg_inf;
  wire p1_data_enable;
  wire p1_not_valid;
  wire [22:0] FRACTION_HIGH_BIT;
  wire [22:0] sign_ext_92833;
  wire [7:0] MAX_EXPONENT__2;
  wire [8:0] add_92774;
  wire [27:0] shrl_92780;
  wire [26:0] shifted_fraction;
  wire [2:0] concat_92663;
  wire [2:0] concat_92664;
  wire [2:0] concat_92665;
  wire [1:0] concat_92668;
  wire [2:0] concat_92674;
  wire result_sign__1;
  wire [27:0] neg_92415;
  wire [27:0] wide_y;
  wire p0_enable;
  wire p0_all_active_inputs_valid;
  wire [8:0] sum;
  wire [22:0] result_fraction__4;
  wire [22:0] result_fraction__3;
  wire [7:0] result_exponent__2;
  wire [8:0] wide_exponent__2;
  wire [9:0] concat_92775;
  wire [22:0] result_fraction;
  wire [2:0] normal_chunk;
  wire [1:0] half_way_chunk;
  wire [23:0] bit_slice_92735;
  wire nor_92676;
  wire leading_zeroes__4_to_5;
  wire [2:0] priority_sel_92678;
  wire [1:0] priority_sel_92679;
  wire [2:0] priority_sel_92680;
  wire or_92681;
  wire result_sign__2;
  wire [27:0] abs_fraction;
  wire not_92500;
  wire result_sign;
  wire xor_92419;
  wire [24:0] wide_x_squeezed;
  wire [24:0] bit_slice_92421;
  wire [27:0] shrl_92422;
  wire sticky;
  wire is_operand_inf;
  wire and_92452;
  wire is_result_nan;
  wire not_92454;
  wire p0_data_enable;
  wire bit_slice_92360;
  wire [22:0] tuple_index_92361;
  wire [22:0] tuple_index_92362;
  wire [7:0] bit_slice_92363;
  wire tuple_index_92364;
  wire tuple_index_92365;
  wire [31:0] __xls_float_ips__result_buf;
  assign xls_float_ips__result_valid_inv = ~__xls_float_ips__result_valid_reg;
  assign xls_float_ips__result_valid_load_en = xls_float_ips__result_rdy | xls_float_ips__result_valid_inv;
  assign xls_float_ips__result_load_en = p7_valid & xls_float_ips__result_valid_load_en;
  assign p8_stage_done = p7_valid & xls_float_ips__result_load_en;
  assign p8_not_valid = ~p7_valid;
  assign p7_enable = p8_stage_done | p8_not_valid;
  assign p7_data_enable = p7_enable & p6_valid;
  assign p7_not_valid = ~p6_valid;
  assign p6_enable = p7_data_enable | p7_not_valid;
  assign p6_data_enable = p6_enable & p5_valid;
  assign p6_not_valid = ~p5_valid;
  assign p5_enable = p6_data_enable | p6_not_valid;
  assign p5_data_enable = p5_enable & p4_valid;
  assign p5_not_valid = ~p4_valid;
  assign p4_enable = p5_data_enable | p5_not_valid;
  assign p4_data_enable = p4_enable & p3_valid;
  assign p4_not_valid = ~p3_valid;
  assign fraction_shift__3 = 3'h4;
  assign p3_enable = p4_data_enable | p4_not_valid;
  assign add_92802 = p5_concat_92775 + 10'h001;
  assign concat_92763 = {1'h0, p4_bit_slice_92735};
  assign carry_bit = p2_abs_fraction[27];
  assign addend_x__1_squeezed = p1_xor_92419 ? p1_bit_slice_92421 : p1_wide_x_squeezed;
  assign a_bexp = p0_bit_slice_92360 ? p0_a_bexp__1 : p0_b_bexp__5;
  assign incremented_sum__1 = p0_bit_slice_92363 + 8'h01;
  assign MAX_EXPONENT = 8'hff;
  assign a_fraction = p0_bit_slice_92360 ? p0_tuple_index_92362 : p0_tuple_index_92361;
  assign b_bexp = p0_bit_slice_92360 ? p0_b_bexp__5 : p0_a_bexp__1;
  assign MAX_EXPONENT__1 = 8'hff;
  assign b_fraction = p0_bit_slice_92360 ? p0_tuple_index_92361 : p0_tuple_index_92362;
  assign p3_data_enable = p3_enable & p2_valid;
  assign p3_not_valid = ~p2_valid;
  assign wide_exponent = add_92802 - {5'h00, p5_leading_zeroes__4_to_5, p5_leading_zeroes__0_to_4};
  assign do_round_up = p4_normal_chunk > fraction_shift__3 | p4_half_way_chunk == 2'h3;
  assign add_92766 = concat_92763 + 25'h000_0001;
  assign leading_zeroes__0_to_4 = priority_sel_4b_2way({p3_nor_92676, p3_leading_zeroes__4_to_5}, {p3_and_92643, p3_priority_sel_92678}, {1'h1, p3_nor_92649, p3_priority_sel_92679}, {p3_and_92641, p3_priority_sel_92680});
  assign nor_92548 = ~(p2_abs_fraction[11] | p2_abs_fraction[10]);
  assign nor_92549 = ~(p2_abs_fraction[9] | p2_abs_fraction[8]);
  assign nor_92551 = ~(p2_abs_fraction[1] | p2_abs_fraction[0]);
  assign nor_92552 = ~(p2_abs_fraction[3] | p2_abs_fraction[2]);
  assign nor_92557 = ~(p2_abs_fraction[5] | p2_abs_fraction[4]);
  assign nor_92558 = ~(p2_abs_fraction[7] | p2_abs_fraction[6]);
  assign nor_92563 = ~(p2_abs_fraction[17] | p2_abs_fraction[16]);
  assign nor_92566 = ~(p2_abs_fraction[13] | p2_abs_fraction[12]);
  assign nor_92567 = ~(carry_bit | p2_abs_fraction[26]);
  assign nor_92568 = ~(p2_abs_fraction[25] | p2_abs_fraction[24]);
  assign nor_92574 = ~(p2_abs_fraction[21] | p2_abs_fraction[20]);
  assign a_bexpbs_difference__1 = p0_bit_slice_92360 ? incremented_sum__1 : ~p0_bit_slice_92363;
  assign eq_92432 = a_bexp == MAX_EXPONENT;
  assign eq_92433 = a_fraction == 23'h00_0000;
  assign eq_92434 = b_bexp == MAX_EXPONENT__1;
  assign eq_92435 = b_fraction == 23'h00_0000;
  assign p2_enable = p3_data_enable | p3_not_valid;
  assign and_reduce_92829 = &p6_wide_exponent__2[7:0];
  assign wide_exponent__1 = wide_exponent & {10{p5_not_92500}};
  assign rounded_fraction_squeezed_portion_3_width_25 = do_round_up ? add_92766 : concat_92763;
  assign leading_zeroes = {p3_leading_zeroes__4_to_5, leading_zeroes__0_to_4};
  assign nor_92575 = ~(p2_abs_fraction[23] | p2_abs_fraction[22]);
  assign and_92576 = nor_92548 & nor_92549;
  assign and_92578 = nor_92552 & nor_92551;
  assign nor_92583 = ~(p2_abs_fraction[7] | p2_abs_fraction[6] | nor_92557);
  assign and_92584 = nor_92558 & nor_92557;
  assign nor_92587 = ~(p2_abs_fraction[11] | ~p2_abs_fraction[10]);
  assign and_92591 = ~(p2_abs_fraction[19] | p2_abs_fraction[18]) & nor_92563;
  assign nor_92592 = ~(p2_abs_fraction[15] | p2_abs_fraction[14]);
  assign and_92596 = nor_92567 & nor_92568;
  assign nor_92598 = ~(carry_bit | ~p2_abs_fraction[26]);
  assign add_92484 = {{1{addend_x__1_squeezed[24]}}, addend_x__1_squeezed} + {1'h0, p1_shrl_92422[27:3]};
  assign fraction_x = {1'h1, a_fraction};
  assign a_sign = p0_bit_slice_92360 ? p0_tuple_index_92365 : p0_tuple_index_92364;
  assign b_sign = p0_bit_slice_92360 ? p0_tuple_index_92364 : p0_tuple_index_92365;
  assign p2_data_enable = p2_enable & p1_valid;
  assign p2_not_valid = ~p1_valid;
  assign b_bexp__5 = xls_float_ips__rhs[30:23];
  assign rounding_carry = rounded_fraction_squeezed_portion_3_width_25[24];
  assign fraction_shift__2 = 3'h3;
  assign fraction_shift__4 = 3'h4;
  assign cancel_fraction = leading_zeroes >= 5'h1d ? 29'h0000_0000 : {1'h0, p3_abs_fraction} << leading_zeroes;
  assign and_92605 = nor_92575 & nor_92574;
  assign and_92623 = nor_92592 & nor_92566;
  assign fraction_x__1 = fraction_x & {24{a_bexp != 8'h00}};
  assign addend_x__1_squeezed_const_lsb_bits__1 = 3'h0;
  assign fraction_y = {1'h1, b_fraction};
  assign sign_ext_92404 = {24{b_bexp != 8'h00}};
  assign add_92423 = (a_bexpbs_difference__1 >= 8'h1c ? 28'h000_0000 : 28'h000_0001 << a_bexpbs_difference__1) + 28'hfff_ffff;
  assign p1_enable = p2_data_enable | p2_not_valid;
  assign a_bexp__1 = xls_float_ips__lhs[30:23];
  assign rounded_fraction = {rounded_fraction_squeezed_portion_3_width_25, p4_normal_chunk};
  assign fraction_shift__1 = rounding_carry ? fraction_shift__4 : fraction_shift__2;
  assign cancel_fraction__1 = cancel_fraction[27:1];
  assign carry_fraction__1 = {p3_abs_fraction[27:2], p3_or_92681};
  assign and_92641 = and_92596 & and_92605;
  assign and_92643 = and_92576 & and_92584;
  assign nor_92649 = ~(~and_92591 | and_92623);
  assign and_92650 = and_92591 & and_92623;
  assign priority_sel_92657 = priority_sel_2b_2way({~(carry_bit | p2_abs_fraction[26] | nor_92568), and_92596}, {nor_92598, 1'h0}, {1'h1, ~(p2_abs_fraction[25] | ~p2_abs_fraction[24])}, {nor_92567, nor_92598});
  assign concat_92489 = {add_92484[24:0], p1_shrl_92422[2:1], p1_shrl_92422[0] | p1_sticky};
  assign fraction_is_zero = add_92484 == 26'h000_0000 & ~(p1_shrl_92422[1] | p1_shrl_92422[2]) & ~(p1_shrl_92422[0] | p1_sticky);
  assign wide_x = {1'h0, fraction_x__1, addend_x__1_squeezed_const_lsb_bits__1};
  assign fraction_y__1 = fraction_y & sign_ext_92404;
  assign addend_x__1_squeezed_const_lsb_bits = 3'h0;
  assign has_pos_inf = ~(~eq_92432 | ~eq_92433 | a_sign) | ~(~eq_92434 | ~eq_92435 | b_sign);
  assign has_neg_inf = eq_92432 & eq_92433 & a_sign | eq_92434 & eq_92435 & b_sign;
  assign p1_data_enable = p1_enable & p0_valid;
  assign p1_not_valid = ~p0_valid;
  assign FRACTION_HIGH_BIT = 23'h40_0000;
  assign sign_ext_92833 = {23{~(p6_is_operand_inf | p6_wide_exponent__2[8] | and_reduce_92829 | ~((|p6_wide_exponent__2[8:1]) | p6_wide_exponent__2[0]))}};
  assign MAX_EXPONENT__2 = 8'hff;
  assign add_92774 = {1'h0, p4_a_bexp} + {8'h00, rounding_carry};
  assign shrl_92780 = rounded_fraction >> fraction_shift__1;
  assign shifted_fraction = p3_carry_bit ? carry_fraction__1 : cancel_fraction__1;
  assign concat_92663 = {and_92578, priority_sel_2b_2way({~(p2_abs_fraction[3] | p2_abs_fraction[2] | nor_92551), and_92578}, 2'h0, {1'h1, ~(p2_abs_fraction[1] | ~p2_abs_fraction[0])}, {nor_92552, ~(p2_abs_fraction[3] | ~p2_abs_fraction[2])})};
  assign concat_92664 = {1'h1, nor_92583, priority_sel_1b_4way({~(p2_abs_fraction[7] | ~p2_abs_fraction[6]), nor_92558, nor_92583, and_92584}, 1'h0, ~(p2_abs_fraction[5] | ~p2_abs_fraction[4]), 1'h0, 1'h1, 1'h0)};
  assign concat_92665 = {and_92576, priority_sel_2b_2way({~(p2_abs_fraction[11] | p2_abs_fraction[10] | nor_92549), and_92576}, {nor_92587, 1'h0}, {1'h1, ~(p2_abs_fraction[9] | ~p2_abs_fraction[8])}, {nor_92548, nor_92587})};
  assign concat_92668 = {nor_92592, priority_sel_1b_3way({~(p2_abs_fraction[15] | ~p2_abs_fraction[14]), nor_92592, ~(p2_abs_fraction[15] | p2_abs_fraction[14] | nor_92566)}, ~(p2_abs_fraction[13] | ~p2_abs_fraction[12]), 1'h0, 1'h1, 1'h0)};
  assign concat_92674 = {1'h1, nor_92575, priority_sel_1b_3way({~(p2_abs_fraction[23] | ~p2_abs_fraction[22]), nor_92575, ~(p2_abs_fraction[23] | p2_abs_fraction[22] | nor_92574)}, ~(p2_abs_fraction[21] | ~p2_abs_fraction[20]), 1'h0, 1'h1, 1'h0)};
  assign result_sign__1 = p2_is_operand_inf ? p2_not_92454 : p2_result_sign;
  assign neg_92415 = -wide_x;
  assign wide_y = {1'h0, fraction_y__1, addend_x__1_squeezed_const_lsb_bits};
  assign p0_enable = p1_data_enable | p1_not_valid;
  assign p0_all_active_inputs_valid = xls_float_ips__rhs_vld & xls_float_ips__lhs_vld;
  assign sum = {1'h0, a_bexp__1} + {1'h0, ~b_bexp__5};
  assign result_fraction__4 = p7_is_result_nan ? FRACTION_HIGH_BIT : p7_result_fraction__3;
  assign result_fraction__3 = p6_result_fraction & sign_ext_92833;
  assign result_exponent__2 = p6_is_result_nan | p6_is_operand_inf | p6_wide_exponent__2[8] | and_reduce_92829 ? MAX_EXPONENT__2 : p6_wide_exponent__2[7:0];
  assign wide_exponent__2 = wide_exponent__1[8:0] & {9{~wide_exponent__1[9]}};
  assign concat_92775 = {1'h0, add_92774};
  assign result_fraction = shrl_92780[22:0];
  assign normal_chunk = shifted_fraction[2:0];
  assign half_way_chunk = shifted_fraction[3:2];
  assign bit_slice_92735 = shifted_fraction[26:3];
  assign nor_92676 = ~(~and_92641 | and_92650);
  assign leading_zeroes__4_to_5 = and_92641 & and_92650;
  assign priority_sel_92678 = priority_sel_3b_2way({~(~and_92576 | and_92584), and_92643}, concat_92663, concat_92664, concat_92665);
  assign priority_sel_92679 = priority_sel_2b_4way({~(p2_abs_fraction[19] | p2_abs_fraction[18] | nor_92563), and_92591, nor_92649, and_92650}, 2'h0, concat_92668, 2'h0, {1'h1, ~(p2_abs_fraction[17] | ~p2_abs_fraction[16])}, {1'h0, ~(p2_abs_fraction[19] | ~p2_abs_fraction[18])});
  assign priority_sel_92680 = priority_sel_3b_2way({~(~and_92596 | and_92605), and_92641}, {priority_sel_92657, 1'h0}, concat_92674, {and_92596, priority_sel_92657});
  assign or_92681 = p2_abs_fraction[1] | p2_abs_fraction[0];
  assign result_sign__2 = ~p2_is_result_nan & result_sign__1;
  assign abs_fraction = add_92484[25] ? -concat_92489 : concat_92489;
  assign not_92500 = ~fraction_is_zero;
  assign result_sign = priority_sel_1b_2way({add_92484[25], fraction_is_zero}, p1_and_92452, ~p1_b_sign, p1_b_sign);
  assign xor_92419 = a_sign ^ b_sign;
  assign wide_x_squeezed = {1'h0, fraction_x__1};
  assign bit_slice_92421 = neg_92415[27:3];
  assign shrl_92422 = a_bexpbs_difference__1 >= 8'h1c ? 28'h000_0000 : wide_y >> a_bexpbs_difference__1;
  assign sticky = (fraction_y & sign_ext_92404 & add_92423[26:3]) != 24'h00_0000;
  assign is_operand_inf = eq_92432 & eq_92433 | eq_92434 & eq_92435;
  assign and_92452 = a_sign & b_sign;
  assign is_result_nan = ~(~eq_92432 | eq_92433) | ~(~eq_92434 | eq_92435) | has_pos_inf & has_neg_inf;
  assign not_92454 = ~has_pos_inf;
  assign p0_data_enable = p0_enable & p0_all_active_inputs_valid;
  assign bit_slice_92360 = sum[8];
  assign tuple_index_92361 = xls_float_ips__rhs[22:0];
  assign tuple_index_92362 = xls_float_ips__lhs[22:0];
  assign bit_slice_92363 = sum[7:0];
  assign tuple_index_92364 = xls_float_ips__rhs[31:31];
  assign tuple_index_92365 = xls_float_ips__lhs[31:31];
  assign __xls_float_ips__result_buf = {p7_result_sign__2, p7_result_exponent__2, result_fraction__4};
  always @ (posedge clk) begin
    if (rst) begin
      p0_b_bexp__5 <= 8'h00;
      p0_a_bexp__1 <= 8'h00;
      p0_bit_slice_92360 <= 1'h0;
      p0_tuple_index_92361 <= 23'h00_0000;
      p0_tuple_index_92362 <= 23'h00_0000;
      p0_bit_slice_92363 <= 8'h00;
      p0_tuple_index_92364 <= 1'h0;
      p0_tuple_index_92365 <= 1'h0;
      p1_a_bexp <= 8'h00;
      p1_b_sign <= 1'h0;
      p1_xor_92419 <= 1'h0;
      p1_wide_x_squeezed <= 25'h000_0000;
      p1_bit_slice_92421 <= 25'h000_0000;
      p1_shrl_92422 <= 28'h000_0000;
      p1_sticky <= 1'h0;
      p1_is_operand_inf <= 1'h0;
      p1_and_92452 <= 1'h0;
      p1_is_result_nan <= 1'h0;
      p1_not_92454 <= 1'h0;
      p2_a_bexp <= 8'h00;
      p2_abs_fraction <= 28'h000_0000;
      p2_not_92500 <= 1'h0;
      p2_is_operand_inf <= 1'h0;
      p2_is_result_nan <= 1'h0;
      p2_result_sign <= 1'h0;
      p2_not_92454 <= 1'h0;
      p3_a_bexp <= 8'h00;
      p3_abs_fraction <= 28'h000_0000;
      p3_carry_bit <= 1'h0;
      p3_and_92641 <= 1'h0;
      p3_and_92643 <= 1'h0;
      p3_nor_92649 <= 1'h0;
      p3_nor_92676 <= 1'h0;
      p3_leading_zeroes__4_to_5 <= 1'h0;
      p3_priority_sel_92678 <= 3'h0;
      p3_priority_sel_92679 <= 2'h0;
      p3_priority_sel_92680 <= 3'h0;
      p3_or_92681 <= 1'h0;
      p3_not_92500 <= 1'h0;
      p3_is_operand_inf <= 1'h0;
      p3_is_result_nan <= 1'h0;
      p3_result_sign__2 <= 1'h0;
      p4_a_bexp <= 8'h00;
      p4_leading_zeroes__4_to_5 <= 1'h0;
      p4_leading_zeroes__0_to_4 <= 4'h0;
      p4_normal_chunk <= 3'h0;
      p4_half_way_chunk <= 2'h0;
      p4_bit_slice_92735 <= 24'h00_0000;
      p4_not_92500 <= 1'h0;
      p4_is_operand_inf <= 1'h0;
      p4_is_result_nan <= 1'h0;
      p4_result_sign__2 <= 1'h0;
      p5_leading_zeroes__4_to_5 <= 1'h0;
      p5_leading_zeroes__0_to_4 <= 4'h0;
      p5_concat_92775 <= 10'h000;
      p5_not_92500 <= 1'h0;
      p5_is_operand_inf <= 1'h0;
      p5_is_result_nan <= 1'h0;
      p5_result_fraction <= 23'h00_0000;
      p5_result_sign__2 <= 1'h0;
      p6_wide_exponent__2 <= 9'h000;
      p6_is_operand_inf <= 1'h0;
      p6_is_result_nan <= 1'h0;
      p6_result_fraction <= 23'h00_0000;
      p6_result_sign__2 <= 1'h0;
      p7_is_result_nan <= 1'h0;
      p7_result_fraction__3 <= 23'h00_0000;
      p7_result_sign__2 <= 1'h0;
      p7_result_exponent__2 <= 8'h00;
      p0_valid <= 1'h0;
      p1_valid <= 1'h0;
      p2_valid <= 1'h0;
      p3_valid <= 1'h0;
      p4_valid <= 1'h0;
      p5_valid <= 1'h0;
      p6_valid <= 1'h0;
      p7_valid <= 1'h0;
      __xls_float_ips__result_reg <= __xls_float_ips__result_reg_init;
      __xls_float_ips__result_valid_reg <= 1'h0;
    end else begin
      p0_b_bexp__5 <= p0_data_enable ? b_bexp__5 : p0_b_bexp__5;
      p0_a_bexp__1 <= p0_data_enable ? a_bexp__1 : p0_a_bexp__1;
      p0_bit_slice_92360 <= p0_data_enable ? bit_slice_92360 : p0_bit_slice_92360;
      p0_tuple_index_92361 <= p0_data_enable ? tuple_index_92361 : p0_tuple_index_92361;
      p0_tuple_index_92362 <= p0_data_enable ? tuple_index_92362 : p0_tuple_index_92362;
      p0_bit_slice_92363 <= p0_data_enable ? bit_slice_92363 : p0_bit_slice_92363;
      p0_tuple_index_92364 <= p0_data_enable ? tuple_index_92364 : p0_tuple_index_92364;
      p0_tuple_index_92365 <= p0_data_enable ? tuple_index_92365 : p0_tuple_index_92365;
      p1_a_bexp <= p1_data_enable ? a_bexp : p1_a_bexp;
      p1_b_sign <= p1_data_enable ? b_sign : p1_b_sign;
      p1_xor_92419 <= p1_data_enable ? xor_92419 : p1_xor_92419;
      p1_wide_x_squeezed <= p1_data_enable ? wide_x_squeezed : p1_wide_x_squeezed;
      p1_bit_slice_92421 <= p1_data_enable ? bit_slice_92421 : p1_bit_slice_92421;
      p1_shrl_92422 <= p1_data_enable ? shrl_92422 : p1_shrl_92422;
      p1_sticky <= p1_data_enable ? sticky : p1_sticky;
      p1_is_operand_inf <= p1_data_enable ? is_operand_inf : p1_is_operand_inf;
      p1_and_92452 <= p1_data_enable ? and_92452 : p1_and_92452;
      p1_is_result_nan <= p1_data_enable ? is_result_nan : p1_is_result_nan;
      p1_not_92454 <= p1_data_enable ? not_92454 : p1_not_92454;
      p2_a_bexp <= p2_data_enable ? p1_a_bexp : p2_a_bexp;
      p2_abs_fraction <= p2_data_enable ? abs_fraction : p2_abs_fraction;
      p2_not_92500 <= p2_data_enable ? not_92500 : p2_not_92500;
      p2_is_operand_inf <= p2_data_enable ? p1_is_operand_inf : p2_is_operand_inf;
      p2_is_result_nan <= p2_data_enable ? p1_is_result_nan : p2_is_result_nan;
      p2_result_sign <= p2_data_enable ? result_sign : p2_result_sign;
      p2_not_92454 <= p2_data_enable ? p1_not_92454 : p2_not_92454;
      p3_a_bexp <= p3_data_enable ? p2_a_bexp : p3_a_bexp;
      p3_abs_fraction <= p3_data_enable ? p2_abs_fraction : p3_abs_fraction;
      p3_carry_bit <= p3_data_enable ? carry_bit : p3_carry_bit;
      p3_and_92641 <= p3_data_enable ? and_92641 : p3_and_92641;
      p3_and_92643 <= p3_data_enable ? and_92643 : p3_and_92643;
      p3_nor_92649 <= p3_data_enable ? nor_92649 : p3_nor_92649;
      p3_nor_92676 <= p3_data_enable ? nor_92676 : p3_nor_92676;
      p3_leading_zeroes__4_to_5 <= p3_data_enable ? leading_zeroes__4_to_5 : p3_leading_zeroes__4_to_5;
      p3_priority_sel_92678 <= p3_data_enable ? priority_sel_92678 : p3_priority_sel_92678;
      p3_priority_sel_92679 <= p3_data_enable ? priority_sel_92679 : p3_priority_sel_92679;
      p3_priority_sel_92680 <= p3_data_enable ? priority_sel_92680 : p3_priority_sel_92680;
      p3_or_92681 <= p3_data_enable ? or_92681 : p3_or_92681;
      p3_not_92500 <= p3_data_enable ? p2_not_92500 : p3_not_92500;
      p3_is_operand_inf <= p3_data_enable ? p2_is_operand_inf : p3_is_operand_inf;
      p3_is_result_nan <= p3_data_enable ? p2_is_result_nan : p3_is_result_nan;
      p3_result_sign__2 <= p3_data_enable ? result_sign__2 : p3_result_sign__2;
      p4_a_bexp <= p4_data_enable ? p3_a_bexp : p4_a_bexp;
      p4_leading_zeroes__4_to_5 <= p4_data_enable ? p3_leading_zeroes__4_to_5 : p4_leading_zeroes__4_to_5;
      p4_leading_zeroes__0_to_4 <= p4_data_enable ? leading_zeroes__0_to_4 : p4_leading_zeroes__0_to_4;
      p4_normal_chunk <= p4_data_enable ? normal_chunk : p4_normal_chunk;
      p4_half_way_chunk <= p4_data_enable ? half_way_chunk : p4_half_way_chunk;
      p4_bit_slice_92735 <= p4_data_enable ? bit_slice_92735 : p4_bit_slice_92735;
      p4_not_92500 <= p4_data_enable ? p3_not_92500 : p4_not_92500;
      p4_is_operand_inf <= p4_data_enable ? p3_is_operand_inf : p4_is_operand_inf;
      p4_is_result_nan <= p4_data_enable ? p3_is_result_nan : p4_is_result_nan;
      p4_result_sign__2 <= p4_data_enable ? p3_result_sign__2 : p4_result_sign__2;
      p5_leading_zeroes__4_to_5 <= p5_data_enable ? p4_leading_zeroes__4_to_5 : p5_leading_zeroes__4_to_5;
      p5_leading_zeroes__0_to_4 <= p5_data_enable ? p4_leading_zeroes__0_to_4 : p5_leading_zeroes__0_to_4;
      p5_concat_92775 <= p5_data_enable ? concat_92775 : p5_concat_92775;
      p5_not_92500 <= p5_data_enable ? p4_not_92500 : p5_not_92500;
      p5_is_operand_inf <= p5_data_enable ? p4_is_operand_inf : p5_is_operand_inf;
      p5_is_result_nan <= p5_data_enable ? p4_is_result_nan : p5_is_result_nan;
      p5_result_fraction <= p5_data_enable ? result_fraction : p5_result_fraction;
      p5_result_sign__2 <= p5_data_enable ? p4_result_sign__2 : p5_result_sign__2;
      p6_wide_exponent__2 <= p6_data_enable ? wide_exponent__2 : p6_wide_exponent__2;
      p6_is_operand_inf <= p6_data_enable ? p5_is_operand_inf : p6_is_operand_inf;
      p6_is_result_nan <= p6_data_enable ? p5_is_result_nan : p6_is_result_nan;
      p6_result_fraction <= p6_data_enable ? p5_result_fraction : p6_result_fraction;
      p6_result_sign__2 <= p6_data_enable ? p5_result_sign__2 : p6_result_sign__2;
      p7_is_result_nan <= p7_data_enable ? p6_is_result_nan : p7_is_result_nan;
      p7_result_fraction__3 <= p7_data_enable ? result_fraction__3 : p7_result_fraction__3;
      p7_result_sign__2 <= p7_data_enable ? p6_result_sign__2 : p7_result_sign__2;
      p7_result_exponent__2 <= p7_data_enable ? result_exponent__2 : p7_result_exponent__2;
      p0_valid <= p0_enable ? p0_all_active_inputs_valid : p0_valid;
      p1_valid <= p1_enable ? p0_valid : p1_valid;
      p2_valid <= p2_enable ? p1_valid : p2_valid;
      p3_valid <= p3_enable ? p2_valid : p3_valid;
      p4_valid <= p4_enable ? p3_valid : p4_valid;
      p5_valid <= p5_enable ? p4_valid : p5_valid;
      p6_valid <= p6_enable ? p5_valid : p6_valid;
      p7_valid <= p7_enable ? p6_valid : p7_valid;
      __xls_float_ips__result_reg <= xls_float_ips__result_load_en ? __xls_float_ips__result_buf : __xls_float_ips__result_reg;
      __xls_float_ips__result_valid_reg <= xls_float_ips__result_valid_load_en ? p7_valid : __xls_float_ips__result_valid_reg;
    end
  end
  assign xls_float_ips__result = __xls_float_ips__result_reg;
  assign xls_float_ips__result_vld = __xls_float_ips__result_valid_reg;
  assign xls_float_ips__rhs_rdy = p0_data_enable;
  assign xls_float_ips__lhs_rdy = p0_data_enable;
endmodule
module __xls_float_ips__cmpf32_OEQ_0_next(
  input wire clk,
  input wire rst,
  input wire [31:0] xls_float_ips__lhs,
  input wire xls_float_ips__lhs_vld,
  input wire [31:0] xls_float_ips__rhs,
  input wire xls_float_ips__rhs_vld,
  input wire xls_float_ips__result_rdy,
  output wire xls_float_ips__result,
  output wire xls_float_ips__result_vld,
  output wire xls_float_ips__lhs_rdy,
  output wire xls_float_ips__rhs_rdy
);
  reg __xls_float_ips__result_reg;
  reg __xls_float_ips__result_valid_reg;
  wire [7:0] a_bexp__1;
  wire [22:0] a_fraction__1;
  wire [7:0] b_bexp;
  wire [22:0] b_fraction;
  wire a_sign__1;
  wire b_sign;
  wire xls_float_ips__result_valid_inv;
  wire p0_all_active_inputs_valid;
  wire xls_float_ips__result_valid_load_en;
  wire xls_float_ips__result_load_en;
  wire p0_stage_done;
  wire __xls_float_ips__result_buf;
  assign a_bexp__1 = xls_float_ips__lhs[30:23];
  assign a_fraction__1 = xls_float_ips__lhs[22:0];
  assign b_bexp = xls_float_ips__rhs[30:23];
  assign b_fraction = xls_float_ips__rhs[22:0];
  assign a_sign__1 = xls_float_ips__lhs[31:31];
  assign b_sign = xls_float_ips__rhs[31:31];
  assign xls_float_ips__result_valid_inv = ~__xls_float_ips__result_valid_reg;
  assign p0_all_active_inputs_valid = xls_float_ips__lhs_vld & xls_float_ips__rhs_vld;
  assign xls_float_ips__result_valid_load_en = xls_float_ips__result_rdy | xls_float_ips__result_valid_inv;
  assign xls_float_ips__result_load_en = p0_all_active_inputs_valid & xls_float_ips__result_valid_load_en;
  assign p0_stage_done = p0_all_active_inputs_valid & xls_float_ips__result_load_en;
  assign __xls_float_ips__result_buf = ~(a_bexp__1 == 8'hff & a_fraction__1 != 23'h00_0000 | b_bexp == 8'hff & b_fraction != 23'h00_0000) & (a_sign__1 == b_sign & a_bexp__1 == b_bexp & a_fraction__1 == b_fraction | a_bexp__1 == 8'h00 & b_bexp == 8'h00);
  always @ (posedge clk) begin
    if (rst) begin
      __xls_float_ips__result_reg <= 1'h0;
      __xls_float_ips__result_valid_reg <= 1'h0;
    end else begin
      __xls_float_ips__result_reg <= xls_float_ips__result_load_en ? __xls_float_ips__result_buf : __xls_float_ips__result_reg;
      __xls_float_ips__result_valid_reg <= xls_float_ips__result_valid_load_en ? p0_all_active_inputs_valid : __xls_float_ips__result_valid_reg;
    end
  end
  assign xls_float_ips__result = __xls_float_ips__result_reg;
  assign xls_float_ips__result_vld = __xls_float_ips__result_valid_reg;
  assign xls_float_ips__lhs_rdy = p0_stage_done;
  assign xls_float_ips__rhs_rdy = p0_stage_done;
endmodule
module __xls_float_ips__cmpf32_OGE_0_next(
  input wire clk,
  input wire rst,
  input wire [31:0] xls_float_ips__lhs,
  input wire xls_float_ips__lhs_vld,
  input wire [31:0] xls_float_ips__rhs,
  input wire xls_float_ips__rhs_vld,
  input wire xls_float_ips__result_rdy,
  output wire xls_float_ips__result,
  output wire xls_float_ips__result_vld,
  output wire xls_float_ips__lhs_rdy,
  output wire xls_float_ips__rhs_rdy
);
  function automatic priority_sel_1b_3way (input reg [2:0] sel, input reg case0, input reg case1, input reg case2, input reg default_value);
    begin
      casez (sel)
        3'b??1: begin
          priority_sel_1b_3way = case0;
        end
        3'b?10: begin
          priority_sel_1b_3way = case1;
        end
        3'b100: begin
          priority_sel_1b_3way = case2;
        end
        3'b000: begin
          priority_sel_1b_3way = default_value;
        end
        default: begin
          // Propagate X
          priority_sel_1b_3way = 1'dx;
        end
      endcase
    end
  endfunction
  reg __xls_float_ips__result_reg;
  reg __xls_float_ips__result_valid_reg;
  wire [7:0] a_bexp__1;
  wire [7:0] b_bexp__2;
  wire eq_747;
  wire eq_748;
  wire [22:0] a_fraction__2;
  wire [22:0] b_fraction__2;
  wire a_sign__2;
  wire b_sign__1;
  wire [22:0] a__1_fraction__5;
  wire [22:0] b__1_fraction__5;
  wire eq_767;
  wire eq_exp;
  wire gt_fraction;
  wire and_771;
  wire and_772;
  wire and_774;
  wire gt_exp;
  wire nor_777;
  wire abs_gt;
  wire and_791;
  wire xls_float_ips__result_valid_inv;
  wire result;
  wire p0_all_active_inputs_valid;
  wire xls_float_ips__result_valid_load_en;
  wire xls_float_ips__result_load_en;
  wire p0_stage_done;
  wire __xls_float_ips__result_buf;
  assign a_bexp__1 = xls_float_ips__lhs[30:23];
  assign b_bexp__2 = xls_float_ips__rhs[30:23];
  assign eq_747 = a_bexp__1 == 8'h00;
  assign eq_748 = b_bexp__2 == 8'h00;
  assign a_fraction__2 = xls_float_ips__lhs[22:0];
  assign b_fraction__2 = xls_float_ips__rhs[22:0];
  assign a_sign__2 = xls_float_ips__lhs[31:31];
  assign b_sign__1 = xls_float_ips__rhs[31:31];
  assign a__1_fraction__5 = a_fraction__2 & {23{~eq_747}};
  assign b__1_fraction__5 = b_fraction__2 & {23{~eq_748}};
  assign eq_767 = a_sign__2 == b_sign__1;
  assign eq_exp = a_bexp__1 == b_bexp__2;
  assign gt_fraction = a__1_fraction__5 > b__1_fraction__5;
  assign and_771 = a_bexp__1 == 8'hff & a_fraction__2 != 23'h00_0000;
  assign and_772 = b_bexp__2 == 8'hff & b_fraction__2 != 23'h00_0000;
  assign and_774 = eq_747 & eq_748;
  assign gt_exp = a_bexp__1 > b_bexp__2;
  assign nor_777 = ~(and_771 | and_772);
  assign abs_gt = gt_exp | eq_exp & gt_fraction;
  assign and_791 = ~abs_gt & ~(nor_777 & (eq_767 & eq_exp & a__1_fraction__5 == b__1_fraction__5 | and_774));
  assign xls_float_ips__result_valid_inv = ~__xls_float_ips__result_valid_reg;
  assign result = priority_sel_1b_3way({~(~a_sign__2 | b_sign__1), ~(a_sign__2 | ~b_sign__1), ~(a_sign__2 | b_sign__1)}, abs_gt, 1'h1, 1'h0, and_791);
  assign p0_all_active_inputs_valid = xls_float_ips__lhs_vld & xls_float_ips__rhs_vld;
  assign xls_float_ips__result_valid_load_en = xls_float_ips__result_rdy | xls_float_ips__result_valid_inv;
  assign xls_float_ips__result_load_en = p0_all_active_inputs_valid & xls_float_ips__result_valid_load_en;
  assign p0_stage_done = p0_all_active_inputs_valid & xls_float_ips__result_load_en;
  assign __xls_float_ips__result_buf = ~(and_771 | and_772 | ~result) | nor_777 & (eq_767 & eq_exp & a_fraction__2 == b_fraction__2 | and_774);
  always @ (posedge clk) begin
    if (rst) begin
      __xls_float_ips__result_reg <= 1'h0;
      __xls_float_ips__result_valid_reg <= 1'h0;
    end else begin
      __xls_float_ips__result_reg <= xls_float_ips__result_load_en ? __xls_float_ips__result_buf : __xls_float_ips__result_reg;
      __xls_float_ips__result_valid_reg <= xls_float_ips__result_valid_load_en ? p0_all_active_inputs_valid : __xls_float_ips__result_valid_reg;
    end
  end
  assign xls_float_ips__result = __xls_float_ips__result_reg;
  assign xls_float_ips__result_vld = __xls_float_ips__result_valid_reg;
  assign xls_float_ips__lhs_rdy = p0_stage_done;
  assign xls_float_ips__rhs_rdy = p0_stage_done;
endmodule
module __xls_float_ips__cmpf32_OGT_0_next(
  input wire clk,
  input wire rst,
  input wire [31:0] xls_float_ips__lhs,
  input wire xls_float_ips__lhs_vld,
  input wire [31:0] xls_float_ips__rhs,
  input wire xls_float_ips__rhs_vld,
  input wire xls_float_ips__result_rdy,
  output wire xls_float_ips__result,
  output wire xls_float_ips__result_vld,
  output wire xls_float_ips__lhs_rdy,
  output wire xls_float_ips__rhs_rdy
);
  function automatic priority_sel_1b_3way (input reg [2:0] sel, input reg case0, input reg case1, input reg case2, input reg default_value);
    begin
      casez (sel)
        3'b??1: begin
          priority_sel_1b_3way = case0;
        end
        3'b?10: begin
          priority_sel_1b_3way = case1;
        end
        3'b100: begin
          priority_sel_1b_3way = case2;
        end
        3'b000: begin
          priority_sel_1b_3way = default_value;
        end
        default: begin
          // Propagate X
          priority_sel_1b_3way = 1'dx;
        end
      endcase
    end
  endfunction
  reg __xls_float_ips__result_reg;
  reg __xls_float_ips__result_valid_reg;
  wire [7:0] a_bexp__2;
  wire [7:0] b_bexp__1;
  wire eq_547;
  wire eq_548;
  wire [22:0] a__1_fraction__1;
  wire [22:0] b__1_fraction__1;
  wire eq_exp;
  wire gt_fraction;
  wire and_568;
  wire and_569;
  wire a_sign__1;
  wire b_sign;
  wire gt_exp;
  wire abs_gt;
  wire xls_float_ips__result_valid_inv;
  wire and_590;
  wire p0_all_active_inputs_valid;
  wire xls_float_ips__result_valid_load_en;
  wire result;
  wire xls_float_ips__result_load_en;
  wire p0_stage_done;
  wire __xls_float_ips__result_buf;
  assign a_bexp__2 = xls_float_ips__lhs[30:23];
  assign b_bexp__1 = xls_float_ips__rhs[30:23];
  assign eq_547 = a_bexp__2 == 8'h00;
  assign eq_548 = b_bexp__1 == 8'h00;
  assign a__1_fraction__1 = xls_float_ips__lhs[22:0] & {23{~eq_547}};
  assign b__1_fraction__1 = xls_float_ips__rhs[22:0] & {23{~eq_548}};
  assign eq_exp = a_bexp__2 == b_bexp__1;
  assign gt_fraction = a__1_fraction__1 > b__1_fraction__1;
  assign and_568 = a_bexp__2 == 8'hff & a__1_fraction__1 != 23'h00_0000;
  assign and_569 = b_bexp__1 == 8'hff & b__1_fraction__1 != 23'h00_0000;
  assign a_sign__1 = xls_float_ips__lhs[31:31];
  assign b_sign = xls_float_ips__rhs[31:31];
  assign gt_exp = a_bexp__2 > b_bexp__1;
  assign abs_gt = gt_exp | eq_exp & gt_fraction;
  assign xls_float_ips__result_valid_inv = ~__xls_float_ips__result_valid_reg;
  assign and_590 = ~abs_gt & ~(~(and_568 | and_569) & (eq_exp & a__1_fraction__1 == b__1_fraction__1 | eq_547 & eq_548));
  assign p0_all_active_inputs_valid = xls_float_ips__lhs_vld & xls_float_ips__rhs_vld;
  assign xls_float_ips__result_valid_load_en = xls_float_ips__result_rdy | xls_float_ips__result_valid_inv;
  assign result = priority_sel_1b_3way({~(~a_sign__1 | b_sign), ~(a_sign__1 | ~b_sign), ~(a_sign__1 | b_sign)}, abs_gt, 1'h1, 1'h0, and_590);
  assign xls_float_ips__result_load_en = p0_all_active_inputs_valid & xls_float_ips__result_valid_load_en;
  assign p0_stage_done = p0_all_active_inputs_valid & xls_float_ips__result_load_en;
  assign __xls_float_ips__result_buf = ~(and_568 | and_569 | ~result);
  always @ (posedge clk) begin
    if (rst) begin
      __xls_float_ips__result_reg <= 1'h0;
      __xls_float_ips__result_valid_reg <= 1'h0;
    end else begin
      __xls_float_ips__result_reg <= xls_float_ips__result_load_en ? __xls_float_ips__result_buf : __xls_float_ips__result_reg;
      __xls_float_ips__result_valid_reg <= xls_float_ips__result_valid_load_en ? p0_all_active_inputs_valid : __xls_float_ips__result_valid_reg;
    end
  end
  assign xls_float_ips__result = __xls_float_ips__result_reg;
  assign xls_float_ips__result_vld = __xls_float_ips__result_valid_reg;
  assign xls_float_ips__lhs_rdy = p0_stage_done;
  assign xls_float_ips__rhs_rdy = p0_stage_done;
endmodule
module __xls_float_ips__cmpf32_OLE_0_next(
  input wire clk,
  input wire rst,
  input wire [31:0] xls_float_ips__lhs,
  input wire xls_float_ips__lhs_vld,
  input wire [31:0] xls_float_ips__rhs,
  input wire xls_float_ips__rhs_vld,
  input wire xls_float_ips__result_rdy,
  output wire xls_float_ips__result,
  output wire xls_float_ips__result_vld,
  output wire xls_float_ips__lhs_rdy,
  output wire xls_float_ips__rhs_rdy
);
  function automatic priority_sel_1b_3way (input reg [2:0] sel, input reg case0, input reg case1, input reg case2, input reg default_value);
    begin
      casez (sel)
        3'b??1: begin
          priority_sel_1b_3way = case0;
        end
        3'b?10: begin
          priority_sel_1b_3way = case1;
        end
        3'b100: begin
          priority_sel_1b_3way = case2;
        end
        3'b000: begin
          priority_sel_1b_3way = default_value;
        end
        default: begin
          // Propagate X
          priority_sel_1b_3way = 1'dx;
        end
      endcase
    end
  endfunction
  reg __xls_float_ips__result_reg;
  reg __xls_float_ips__result_valid_reg;
  wire [7:0] a_bexp__4;
  wire [7:0] b_bexp__2;
  wire eq_710;
  wire eq_711;
  wire [22:0] a_fraction__1;
  wire [22:0] b_fraction;
  wire [22:0] a__1_fraction__5;
  wire [22:0] b__1_fraction__5;
  wire eq_exp;
  wire gt_fraction;
  wire and_731;
  wire and_732;
  wire a_sign__2;
  wire b_sign__1;
  wire gt_exp;
  wire abs_gt;
  wire and_753;
  wire xls_float_ips__result_valid_inv;
  wire result;
  wire p0_all_active_inputs_valid;
  wire xls_float_ips__result_valid_load_en;
  wire xls_float_ips__result_load_en;
  wire p0_stage_done;
  wire __xls_float_ips__result_buf;
  assign a_bexp__4 = xls_float_ips__lhs[30:23];
  assign b_bexp__2 = xls_float_ips__rhs[30:23];
  assign eq_710 = a_bexp__4 == 8'h00;
  assign eq_711 = b_bexp__2 == 8'h00;
  assign a_fraction__1 = xls_float_ips__lhs[22:0];
  assign b_fraction = xls_float_ips__rhs[22:0];
  assign a__1_fraction__5 = a_fraction__1 & {23{~eq_710}};
  assign b__1_fraction__5 = b_fraction & {23{~eq_711}};
  assign eq_exp = a_bexp__4 == b_bexp__2;
  assign gt_fraction = a__1_fraction__5 > b__1_fraction__5;
  assign and_731 = a_bexp__4 == 8'hff & a_fraction__1 != 23'h00_0000;
  assign and_732 = b_bexp__2 == 8'hff & b_fraction != 23'h00_0000;
  assign a_sign__2 = xls_float_ips__lhs[31:31];
  assign b_sign__1 = xls_float_ips__rhs[31:31];
  assign gt_exp = a_bexp__4 > b_bexp__2;
  assign abs_gt = gt_exp | eq_exp & gt_fraction;
  assign and_753 = ~abs_gt & ~(~(and_731 | and_732) & (eq_exp & a__1_fraction__5 == b__1_fraction__5 | eq_710 & eq_711));
  assign xls_float_ips__result_valid_inv = ~__xls_float_ips__result_valid_reg;
  assign result = priority_sel_1b_3way({~(~a_sign__2 | b_sign__1), ~(a_sign__2 | ~b_sign__1), ~(a_sign__2 | b_sign__1)}, abs_gt, 1'h1, 1'h0, and_753);
  assign p0_all_active_inputs_valid = xls_float_ips__lhs_vld & xls_float_ips__rhs_vld;
  assign xls_float_ips__result_valid_load_en = xls_float_ips__result_rdy | xls_float_ips__result_valid_inv;
  assign xls_float_ips__result_load_en = p0_all_active_inputs_valid & xls_float_ips__result_valid_load_en;
  assign p0_stage_done = p0_all_active_inputs_valid & xls_float_ips__result_load_en;
  assign __xls_float_ips__result_buf = ~(and_731 | and_732 | ~(and_731 | and_732 | ~result));
  always @ (posedge clk) begin
    if (rst) begin
      __xls_float_ips__result_reg <= 1'h0;
      __xls_float_ips__result_valid_reg <= 1'h0;
    end else begin
      __xls_float_ips__result_reg <= xls_float_ips__result_load_en ? __xls_float_ips__result_buf : __xls_float_ips__result_reg;
      __xls_float_ips__result_valid_reg <= xls_float_ips__result_valid_load_en ? p0_all_active_inputs_valid : __xls_float_ips__result_valid_reg;
    end
  end
  assign xls_float_ips__result = __xls_float_ips__result_reg;
  assign xls_float_ips__result_vld = __xls_float_ips__result_valid_reg;
  assign xls_float_ips__lhs_rdy = p0_stage_done;
  assign xls_float_ips__rhs_rdy = p0_stage_done;
endmodule
module __xls_float_ips__cmpf32_OLT_0_next(
  input wire clk,
  input wire rst,
  input wire [31:0] xls_float_ips__lhs,
  input wire xls_float_ips__lhs_vld,
  input wire [31:0] xls_float_ips__rhs,
  input wire xls_float_ips__rhs_vld,
  input wire xls_float_ips__result_rdy,
  output wire xls_float_ips__result,
  output wire xls_float_ips__result_vld,
  output wire xls_float_ips__lhs_rdy,
  output wire xls_float_ips__rhs_rdy
);
  function automatic priority_sel_1b_3way (input reg [2:0] sel, input reg case0, input reg case1, input reg case2, input reg default_value);
    begin
      casez (sel)
        3'b??1: begin
          priority_sel_1b_3way = case0;
        end
        3'b?10: begin
          priority_sel_1b_3way = case1;
        end
        3'b100: begin
          priority_sel_1b_3way = case2;
        end
        3'b000: begin
          priority_sel_1b_3way = default_value;
        end
        default: begin
          // Propagate X
          priority_sel_1b_3way = 1'dx;
        end
      endcase
    end
  endfunction
  reg __xls_float_ips__result_reg;
  reg __xls_float_ips__result_valid_reg;
  wire [7:0] a_bexp__4;
  wire [7:0] b_bexp__1;
  wire eq_946;
  wire eq_947;
  wire [22:0] a_fraction__5;
  wire [22:0] b_fraction__1;
  wire a_sign__1;
  wire b_sign__2;
  wire [22:0] a__1_fraction__1;
  wire [22:0] b__1_fraction__1;
  wire eq_966;
  wire eq_exp;
  wire gt_fraction;
  wire and_970;
  wire and_971;
  wire and_973;
  wire gt_exp;
  wire nor_976;
  wire abs_gt;
  wire and_990;
  wire result;
  wire xls_float_ips__result_valid_inv;
  wire p0_all_active_inputs_valid;
  wire xls_float_ips__result_valid_load_en;
  wire xls_float_ips__result_load_en;
  wire p0_stage_done;
  wire __xls_float_ips__result_buf;
  assign a_bexp__4 = xls_float_ips__lhs[30:23];
  assign b_bexp__1 = xls_float_ips__rhs[30:23];
  assign eq_946 = a_bexp__4 == 8'h00;
  assign eq_947 = b_bexp__1 == 8'h00;
  assign a_fraction__5 = xls_float_ips__lhs[22:0];
  assign b_fraction__1 = xls_float_ips__rhs[22:0];
  assign a_sign__1 = xls_float_ips__lhs[31:31];
  assign b_sign__2 = xls_float_ips__rhs[31:31];
  assign a__1_fraction__1 = a_fraction__5 & {23{~eq_946}};
  assign b__1_fraction__1 = b_fraction__1 & {23{~eq_947}};
  assign eq_966 = a_sign__1 == b_sign__2;
  assign eq_exp = a_bexp__4 == b_bexp__1;
  assign gt_fraction = a__1_fraction__1 > b__1_fraction__1;
  assign and_970 = a_bexp__4 == 8'hff & a_fraction__5 != 23'h00_0000;
  assign and_971 = b_bexp__1 == 8'hff & b_fraction__1 != 23'h00_0000;
  assign and_973 = eq_946 & eq_947;
  assign gt_exp = a_bexp__4 > b_bexp__1;
  assign nor_976 = ~(and_970 | and_971);
  assign abs_gt = gt_exp | eq_exp & gt_fraction;
  assign and_990 = ~abs_gt & ~(nor_976 & (eq_966 & eq_exp & a__1_fraction__1 == b__1_fraction__1 | and_973));
  assign result = priority_sel_1b_3way({~(~a_sign__1 | b_sign__2), ~(a_sign__1 | ~b_sign__2), ~(a_sign__1 | b_sign__2)}, abs_gt, 1'h1, 1'h0, and_990);
  assign xls_float_ips__result_valid_inv = ~__xls_float_ips__result_valid_reg;
  assign p0_all_active_inputs_valid = xls_float_ips__lhs_vld & xls_float_ips__rhs_vld;
  assign xls_float_ips__result_valid_load_en = xls_float_ips__result_rdy | xls_float_ips__result_valid_inv;
  assign xls_float_ips__result_load_en = p0_all_active_inputs_valid & xls_float_ips__result_valid_load_en;
  assign p0_stage_done = p0_all_active_inputs_valid & xls_float_ips__result_load_en;
  assign __xls_float_ips__result_buf = ~(and_970 | and_971 | (~(and_970 | and_971 | ~result) | nor_976 & (eq_966 & eq_exp & a_fraction__5 == b_fraction__1 | and_973)));
  always @ (posedge clk) begin
    if (rst) begin
      __xls_float_ips__result_reg <= 1'h0;
      __xls_float_ips__result_valid_reg <= 1'h0;
    end else begin
      __xls_float_ips__result_reg <= xls_float_ips__result_load_en ? __xls_float_ips__result_buf : __xls_float_ips__result_reg;
      __xls_float_ips__result_valid_reg <= xls_float_ips__result_valid_load_en ? p0_all_active_inputs_valid : __xls_float_ips__result_valid_reg;
    end
  end
  assign xls_float_ips__result = __xls_float_ips__result_reg;
  assign xls_float_ips__result_vld = __xls_float_ips__result_valid_reg;
  assign xls_float_ips__lhs_rdy = p0_stage_done;
  assign xls_float_ips__rhs_rdy = p0_stage_done;
endmodule
module __xls_float_ips__cmpf32_UEQ_0_next(
  input wire clk,
  input wire rst,
  input wire [31:0] xls_float_ips__lhs,
  input wire xls_float_ips__lhs_vld,
  input wire [31:0] xls_float_ips__rhs,
  input wire xls_float_ips__rhs_vld,
  input wire xls_float_ips__result_rdy,
  output wire xls_float_ips__result,
  output wire xls_float_ips__result_vld,
  output wire xls_float_ips__lhs_rdy,
  output wire xls_float_ips__rhs_rdy
);
  reg __xls_float_ips__result_reg;
  reg __xls_float_ips__result_valid_reg;
  wire [7:0] a_bexp__1;
  wire [22:0] a_fraction__1;
  wire [7:0] b_bexp__1;
  wire [22:0] b_fraction__1;
  wire a_sign__1;
  wire b_sign;
  wire xls_float_ips__result_valid_inv;
  wire and_265;
  wire and_266;
  wire p0_all_active_inputs_valid;
  wire xls_float_ips__result_valid_load_en;
  wire xls_float_ips__result_load_en;
  wire p0_stage_done;
  wire __xls_float_ips__result_buf;
  assign a_bexp__1 = xls_float_ips__lhs[30:23];
  assign a_fraction__1 = xls_float_ips__lhs[22:0];
  assign b_bexp__1 = xls_float_ips__rhs[30:23];
  assign b_fraction__1 = xls_float_ips__rhs[22:0];
  assign a_sign__1 = xls_float_ips__lhs[31:31];
  assign b_sign = xls_float_ips__rhs[31:31];
  assign xls_float_ips__result_valid_inv = ~__xls_float_ips__result_valid_reg;
  assign and_265 = a_bexp__1 == 8'hff & a_fraction__1 != 23'h00_0000;
  assign and_266 = b_bexp__1 == 8'hff & b_fraction__1 != 23'h00_0000;
  assign p0_all_active_inputs_valid = xls_float_ips__lhs_vld & xls_float_ips__rhs_vld;
  assign xls_float_ips__result_valid_load_en = xls_float_ips__result_rdy | xls_float_ips__result_valid_inv;
  assign xls_float_ips__result_load_en = p0_all_active_inputs_valid & xls_float_ips__result_valid_load_en;
  assign p0_stage_done = p0_all_active_inputs_valid & xls_float_ips__result_load_en;
  assign __xls_float_ips__result_buf = and_265 | and_266 | ~(and_265 | and_266) & (a_sign__1 == b_sign & a_bexp__1 == b_bexp__1 & a_fraction__1 == b_fraction__1 | a_bexp__1 == 8'h00 & b_bexp__1 == 8'h00);
  always @ (posedge clk) begin
    if (rst) begin
      __xls_float_ips__result_reg <= 1'h0;
      __xls_float_ips__result_valid_reg <= 1'h0;
    end else begin
      __xls_float_ips__result_reg <= xls_float_ips__result_load_en ? __xls_float_ips__result_buf : __xls_float_ips__result_reg;
      __xls_float_ips__result_valid_reg <= xls_float_ips__result_valid_load_en ? p0_all_active_inputs_valid : __xls_float_ips__result_valid_reg;
    end
  end
  assign xls_float_ips__result = __xls_float_ips__result_reg;
  assign xls_float_ips__result_vld = __xls_float_ips__result_valid_reg;
  assign xls_float_ips__lhs_rdy = p0_stage_done;
  assign xls_float_ips__rhs_rdy = p0_stage_done;
endmodule
module __xls_float_ips__cmpf32_UGE_0_next(
  input wire clk,
  input wire rst,
  input wire [31:0] xls_float_ips__lhs,
  input wire xls_float_ips__lhs_vld,
  input wire [31:0] xls_float_ips__rhs,
  input wire xls_float_ips__rhs_vld,
  input wire xls_float_ips__result_rdy,
  output wire xls_float_ips__result,
  output wire xls_float_ips__result_vld,
  output wire xls_float_ips__lhs_rdy,
  output wire xls_float_ips__rhs_rdy
);
  function automatic priority_sel_1b_3way (input reg [2:0] sel, input reg case0, input reg case1, input reg case2, input reg default_value);
    begin
      casez (sel)
        3'b??1: begin
          priority_sel_1b_3way = case0;
        end
        3'b?10: begin
          priority_sel_1b_3way = case1;
        end
        3'b100: begin
          priority_sel_1b_3way = case2;
        end
        3'b000: begin
          priority_sel_1b_3way = default_value;
        end
        default: begin
          // Propagate X
          priority_sel_1b_3way = 1'dx;
        end
      endcase
    end
  endfunction
  reg __xls_float_ips__result_reg;
  reg __xls_float_ips__result_valid_reg;
  wire [7:0] a_bexp__1;
  wire [7:0] b_bexp__2;
  wire eq_784;
  wire eq_785;
  wire [22:0] a_fraction__2;
  wire [22:0] b_fraction__2;
  wire a_sign__2;
  wire b_sign__1;
  wire [22:0] a__1_fraction__5;
  wire [22:0] b__1_fraction__5;
  wire eq_804;
  wire eq_exp;
  wire gt_fraction;
  wire and_808;
  wire and_809;
  wire and_811;
  wire gt_exp;
  wire nor_814;
  wire abs_gt;
  wire and_828;
  wire result;
  wire xls_float_ips__result_valid_inv;
  wire p0_all_active_inputs_valid;
  wire xls_float_ips__result_valid_load_en;
  wire not_837;
  wire xls_float_ips__result_load_en;
  wire p0_stage_done;
  wire __xls_float_ips__result_buf;
  assign a_bexp__1 = xls_float_ips__lhs[30:23];
  assign b_bexp__2 = xls_float_ips__rhs[30:23];
  assign eq_784 = a_bexp__1 == 8'h00;
  assign eq_785 = b_bexp__2 == 8'h00;
  assign a_fraction__2 = xls_float_ips__lhs[22:0];
  assign b_fraction__2 = xls_float_ips__rhs[22:0];
  assign a_sign__2 = xls_float_ips__lhs[31:31];
  assign b_sign__1 = xls_float_ips__rhs[31:31];
  assign a__1_fraction__5 = a_fraction__2 & {23{~eq_784}};
  assign b__1_fraction__5 = b_fraction__2 & {23{~eq_785}};
  assign eq_804 = a_sign__2 == b_sign__1;
  assign eq_exp = a_bexp__1 == b_bexp__2;
  assign gt_fraction = a__1_fraction__5 > b__1_fraction__5;
  assign and_808 = a_bexp__1 == 8'hff & a_fraction__2 != 23'h00_0000;
  assign and_809 = b_bexp__2 == 8'hff & b_fraction__2 != 23'h00_0000;
  assign and_811 = eq_784 & eq_785;
  assign gt_exp = a_bexp__1 > b_bexp__2;
  assign nor_814 = ~(and_808 | and_809);
  assign abs_gt = gt_exp | eq_exp & gt_fraction;
  assign and_828 = ~abs_gt & ~(nor_814 & (eq_804 & eq_exp & a__1_fraction__5 == b__1_fraction__5 | and_811));
  assign result = priority_sel_1b_3way({~(~a_sign__2 | b_sign__1), ~(a_sign__2 | ~b_sign__1), ~(a_sign__2 | b_sign__1)}, abs_gt, 1'h1, 1'h0, and_828);
  assign xls_float_ips__result_valid_inv = ~__xls_float_ips__result_valid_reg;
  assign p0_all_active_inputs_valid = xls_float_ips__lhs_vld & xls_float_ips__rhs_vld;
  assign xls_float_ips__result_valid_load_en = xls_float_ips__result_rdy | xls_float_ips__result_valid_inv;
  assign not_837 = ~(~(and_808 | and_809 | ~result) | nor_814 & (eq_804 & eq_exp & a_fraction__2 == b_fraction__2 | and_811));
  assign xls_float_ips__result_load_en = p0_all_active_inputs_valid & xls_float_ips__result_valid_load_en;
  assign p0_stage_done = p0_all_active_inputs_valid & xls_float_ips__result_load_en;
  assign __xls_float_ips__result_buf = and_808 | and_809 | ~(and_808 | and_809 | not_837);
  always @ (posedge clk) begin
    if (rst) begin
      __xls_float_ips__result_reg <= 1'h0;
      __xls_float_ips__result_valid_reg <= 1'h0;
    end else begin
      __xls_float_ips__result_reg <= xls_float_ips__result_load_en ? __xls_float_ips__result_buf : __xls_float_ips__result_reg;
      __xls_float_ips__result_valid_reg <= xls_float_ips__result_valid_load_en ? p0_all_active_inputs_valid : __xls_float_ips__result_valid_reg;
    end
  end
  assign xls_float_ips__result = __xls_float_ips__result_reg;
  assign xls_float_ips__result_vld = __xls_float_ips__result_valid_reg;
  assign xls_float_ips__lhs_rdy = p0_stage_done;
  assign xls_float_ips__rhs_rdy = p0_stage_done;
endmodule
module __xls_float_ips__cmpf32_UGT_0_next(
  input wire clk,
  input wire rst,
  input wire [31:0] xls_float_ips__lhs,
  input wire xls_float_ips__lhs_vld,
  input wire [31:0] xls_float_ips__rhs,
  input wire xls_float_ips__rhs_vld,
  input wire xls_float_ips__result_rdy,
  output wire xls_float_ips__result,
  output wire xls_float_ips__result_vld,
  output wire xls_float_ips__lhs_rdy,
  output wire xls_float_ips__rhs_rdy
);
  function automatic priority_sel_1b_3way (input reg [2:0] sel, input reg case0, input reg case1, input reg case2, input reg default_value);
    begin
      casez (sel)
        3'b??1: begin
          priority_sel_1b_3way = case0;
        end
        3'b?10: begin
          priority_sel_1b_3way = case1;
        end
        3'b100: begin
          priority_sel_1b_3way = case2;
        end
        3'b000: begin
          priority_sel_1b_3way = default_value;
        end
        default: begin
          // Propagate X
          priority_sel_1b_3way = 1'dx;
        end
      endcase
    end
  endfunction
  reg __xls_float_ips__result_reg;
  reg __xls_float_ips__result_valid_reg;
  wire [7:0] a_bexp__2;
  wire [7:0] b_bexp__1;
  wire eq_584;
  wire eq_585;
  wire [22:0] a_fraction;
  wire [22:0] b_fraction;
  wire [22:0] a__1_fraction__1;
  wire [22:0] b__1_fraction__1;
  wire eq_exp;
  wire gt_fraction;
  wire and_605;
  wire and_606;
  wire a_sign__1;
  wire b_sign;
  wire gt_exp;
  wire abs_gt;
  wire and_627;
  wire result;
  wire xls_float_ips__result_valid_inv;
  wire p0_all_active_inputs_valid;
  wire xls_float_ips__result_valid_load_en;
  wire xls_float_ips__result_load_en;
  wire p0_stage_done;
  wire __xls_float_ips__result_buf;
  assign a_bexp__2 = xls_float_ips__lhs[30:23];
  assign b_bexp__1 = xls_float_ips__rhs[30:23];
  assign eq_584 = a_bexp__2 == 8'h00;
  assign eq_585 = b_bexp__1 == 8'h00;
  assign a_fraction = xls_float_ips__lhs[22:0];
  assign b_fraction = xls_float_ips__rhs[22:0];
  assign a__1_fraction__1 = a_fraction & {23{~eq_584}};
  assign b__1_fraction__1 = b_fraction & {23{~eq_585}};
  assign eq_exp = a_bexp__2 == b_bexp__1;
  assign gt_fraction = a__1_fraction__1 > b__1_fraction__1;
  assign and_605 = a_bexp__2 == 8'hff & a_fraction != 23'h00_0000;
  assign and_606 = b_bexp__1 == 8'hff & b_fraction != 23'h00_0000;
  assign a_sign__1 = xls_float_ips__lhs[31:31];
  assign b_sign = xls_float_ips__rhs[31:31];
  assign gt_exp = a_bexp__2 > b_bexp__1;
  assign abs_gt = gt_exp | eq_exp & gt_fraction;
  assign and_627 = ~abs_gt & ~(~(and_605 | and_606) & (eq_exp & a__1_fraction__1 == b__1_fraction__1 | eq_584 & eq_585));
  assign result = priority_sel_1b_3way({~(~a_sign__1 | b_sign), ~(a_sign__1 | ~b_sign), ~(a_sign__1 | b_sign)}, abs_gt, 1'h1, 1'h0, and_627);
  assign xls_float_ips__result_valid_inv = ~__xls_float_ips__result_valid_reg;
  assign p0_all_active_inputs_valid = xls_float_ips__lhs_vld & xls_float_ips__rhs_vld;
  assign xls_float_ips__result_valid_load_en = xls_float_ips__result_rdy | xls_float_ips__result_valid_inv;
  assign xls_float_ips__result_load_en = p0_all_active_inputs_valid & xls_float_ips__result_valid_load_en;
  assign p0_stage_done = p0_all_active_inputs_valid & xls_float_ips__result_load_en;
  assign __xls_float_ips__result_buf = and_605 | and_606 | ~(and_605 | and_606 | ~(~(and_605 | and_606 | ~result)));
  always @ (posedge clk) begin
    if (rst) begin
      __xls_float_ips__result_reg <= 1'h0;
      __xls_float_ips__result_valid_reg <= 1'h0;
    end else begin
      __xls_float_ips__result_reg <= xls_float_ips__result_load_en ? __xls_float_ips__result_buf : __xls_float_ips__result_reg;
      __xls_float_ips__result_valid_reg <= xls_float_ips__result_valid_load_en ? p0_all_active_inputs_valid : __xls_float_ips__result_valid_reg;
    end
  end
  assign xls_float_ips__result = __xls_float_ips__result_reg;
  assign xls_float_ips__result_vld = __xls_float_ips__result_valid_reg;
  assign xls_float_ips__lhs_rdy = p0_stage_done;
  assign xls_float_ips__rhs_rdy = p0_stage_done;
endmodule
module __xls_float_ips__cmpf32_ULE_0_next(
  input wire clk,
  input wire rst,
  input wire [31:0] xls_float_ips__lhs,
  input wire xls_float_ips__lhs_vld,
  input wire [31:0] xls_float_ips__rhs,
  input wire xls_float_ips__rhs_vld,
  input wire xls_float_ips__result_rdy,
  output wire xls_float_ips__result,
  output wire xls_float_ips__result_vld,
  output wire xls_float_ips__lhs_rdy,
  output wire xls_float_ips__rhs_rdy
);
  function automatic priority_sel_1b_3way (input reg [2:0] sel, input reg case0, input reg case1, input reg case2, input reg default_value);
    begin
      casez (sel)
        3'b??1: begin
          priority_sel_1b_3way = case0;
        end
        3'b?10: begin
          priority_sel_1b_3way = case1;
        end
        3'b100: begin
          priority_sel_1b_3way = case2;
        end
        3'b000: begin
          priority_sel_1b_3way = default_value;
        end
        default: begin
          // Propagate X
          priority_sel_1b_3way = 1'dx;
        end
      endcase
    end
  endfunction
  reg __xls_float_ips__result_reg;
  reg __xls_float_ips__result_valid_reg;
  wire [7:0] a_bexp__4;
  wire [7:0] b_bexp__2;
  wire eq_746;
  wire eq_747;
  wire [22:0] a_fraction;
  wire [22:0] b_fraction;
  wire [22:0] a__1_fraction__5;
  wire [22:0] b__1_fraction__5;
  wire eq_exp;
  wire gt_fraction;
  wire and_767;
  wire and_768;
  wire a_sign__2;
  wire b_sign__1;
  wire gt_exp;
  wire abs_gt;
  wire and_789;
  wire result;
  wire xls_float_ips__result_valid_inv;
  wire p0_all_active_inputs_valid;
  wire xls_float_ips__result_valid_load_en;
  wire xls_float_ips__result_load_en;
  wire p0_stage_done;
  wire __xls_float_ips__result_buf;
  assign a_bexp__4 = xls_float_ips__lhs[30:23];
  assign b_bexp__2 = xls_float_ips__rhs[30:23];
  assign eq_746 = a_bexp__4 == 8'h00;
  assign eq_747 = b_bexp__2 == 8'h00;
  assign a_fraction = xls_float_ips__lhs[22:0];
  assign b_fraction = xls_float_ips__rhs[22:0];
  assign a__1_fraction__5 = a_fraction & {23{~eq_746}};
  assign b__1_fraction__5 = b_fraction & {23{~eq_747}};
  assign eq_exp = a_bexp__4 == b_bexp__2;
  assign gt_fraction = a__1_fraction__5 > b__1_fraction__5;
  assign and_767 = a_bexp__4 == 8'hff & a_fraction != 23'h00_0000;
  assign and_768 = b_bexp__2 == 8'hff & b_fraction != 23'h00_0000;
  assign a_sign__2 = xls_float_ips__lhs[31:31];
  assign b_sign__1 = xls_float_ips__rhs[31:31];
  assign gt_exp = a_bexp__4 > b_bexp__2;
  assign abs_gt = gt_exp | eq_exp & gt_fraction;
  assign and_789 = ~abs_gt & ~(~(and_767 | and_768) & (eq_exp & a__1_fraction__5 == b__1_fraction__5 | eq_746 & eq_747));
  assign result = priority_sel_1b_3way({~(~a_sign__2 | b_sign__1), ~(a_sign__2 | ~b_sign__1), ~(a_sign__2 | b_sign__1)}, abs_gt, 1'h1, 1'h0, and_789);
  assign xls_float_ips__result_valid_inv = ~__xls_float_ips__result_valid_reg;
  assign p0_all_active_inputs_valid = xls_float_ips__lhs_vld & xls_float_ips__rhs_vld;
  assign xls_float_ips__result_valid_load_en = xls_float_ips__result_rdy | xls_float_ips__result_valid_inv;
  assign xls_float_ips__result_load_en = p0_all_active_inputs_valid & xls_float_ips__result_valid_load_en;
  assign p0_stage_done = p0_all_active_inputs_valid & xls_float_ips__result_load_en;
  assign __xls_float_ips__result_buf = and_767 | and_768 | ~(and_767 | and_768 | ~(and_767 | and_768 | ~result));
  always @ (posedge clk) begin
    if (rst) begin
      __xls_float_ips__result_reg <= 1'h0;
      __xls_float_ips__result_valid_reg <= 1'h0;
    end else begin
      __xls_float_ips__result_reg <= xls_float_ips__result_load_en ? __xls_float_ips__result_buf : __xls_float_ips__result_reg;
      __xls_float_ips__result_valid_reg <= xls_float_ips__result_valid_load_en ? p0_all_active_inputs_valid : __xls_float_ips__result_valid_reg;
    end
  end
  assign xls_float_ips__result = __xls_float_ips__result_reg;
  assign xls_float_ips__result_vld = __xls_float_ips__result_valid_reg;
  assign xls_float_ips__lhs_rdy = p0_stage_done;
  assign xls_float_ips__rhs_rdy = p0_stage_done;
endmodule
module __xls_float_ips__cmpf32_ULT_0_next(
  input wire clk,
  input wire rst,
  input wire [31:0] xls_float_ips__lhs,
  input wire xls_float_ips__lhs_vld,
  input wire [31:0] xls_float_ips__rhs,
  input wire xls_float_ips__rhs_vld,
  input wire xls_float_ips__result_rdy,
  output wire xls_float_ips__result,
  output wire xls_float_ips__result_vld,
  output wire xls_float_ips__lhs_rdy,
  output wire xls_float_ips__rhs_rdy
);
  function automatic priority_sel_1b_3way (input reg [2:0] sel, input reg case0, input reg case1, input reg case2, input reg default_value);
    begin
      casez (sel)
        3'b??1: begin
          priority_sel_1b_3way = case0;
        end
        3'b?10: begin
          priority_sel_1b_3way = case1;
        end
        3'b100: begin
          priority_sel_1b_3way = case2;
        end
        3'b000: begin
          priority_sel_1b_3way = default_value;
        end
        default: begin
          // Propagate X
          priority_sel_1b_3way = 1'dx;
        end
      endcase
    end
  endfunction
  reg __xls_float_ips__result_reg;
  reg __xls_float_ips__result_valid_reg;
  wire [7:0] a_bexp__4;
  wire [7:0] b_bexp__2;
  wire eq_982;
  wire eq_983;
  wire [22:0] a_fraction__5;
  wire [22:0] b_fraction__2;
  wire a_sign__1;
  wire b_sign__2;
  wire [22:0] a__1_fraction__1;
  wire [22:0] b__1_fraction__1;
  wire eq_1002;
  wire eq_exp;
  wire gt_fraction;
  wire and_1006;
  wire and_1007;
  wire and_1009;
  wire gt_exp;
  wire nor_1012;
  wire abs_gt;
  wire and_1026;
  wire result;
  wire xls_float_ips__result_valid_inv;
  wire p0_all_active_inputs_valid;
  wire xls_float_ips__result_valid_load_en;
  wire xls_float_ips__result_load_en;
  wire nor_1037;
  wire p0_stage_done;
  wire __xls_float_ips__result_buf;
  assign a_bexp__4 = xls_float_ips__lhs[30:23];
  assign b_bexp__2 = xls_float_ips__rhs[30:23];
  assign eq_982 = a_bexp__4 == 8'h00;
  assign eq_983 = b_bexp__2 == 8'h00;
  assign a_fraction__5 = xls_float_ips__lhs[22:0];
  assign b_fraction__2 = xls_float_ips__rhs[22:0];
  assign a_sign__1 = xls_float_ips__lhs[31:31];
  assign b_sign__2 = xls_float_ips__rhs[31:31];
  assign a__1_fraction__1 = a_fraction__5 & {23{~eq_982}};
  assign b__1_fraction__1 = b_fraction__2 & {23{~eq_983}};
  assign eq_1002 = a_sign__1 == b_sign__2;
  assign eq_exp = a_bexp__4 == b_bexp__2;
  assign gt_fraction = a__1_fraction__1 > b__1_fraction__1;
  assign and_1006 = a_bexp__4 == 8'hff & a_fraction__5 != 23'h00_0000;
  assign and_1007 = b_bexp__2 == 8'hff & b_fraction__2 != 23'h00_0000;
  assign and_1009 = eq_982 & eq_983;
  assign gt_exp = a_bexp__4 > b_bexp__2;
  assign nor_1012 = ~(and_1006 | and_1007);
  assign abs_gt = gt_exp | eq_exp & gt_fraction;
  assign and_1026 = ~abs_gt & ~(nor_1012 & (eq_1002 & eq_exp & a__1_fraction__1 == b__1_fraction__1 | and_1009));
  assign result = priority_sel_1b_3way({~(~a_sign__1 | b_sign__2), ~(a_sign__1 | ~b_sign__2), ~(a_sign__1 | b_sign__2)}, abs_gt, 1'h1, 1'h0, and_1026);
  assign xls_float_ips__result_valid_inv = ~__xls_float_ips__result_valid_reg;
  assign p0_all_active_inputs_valid = xls_float_ips__lhs_vld & xls_float_ips__rhs_vld;
  assign xls_float_ips__result_valid_load_en = xls_float_ips__result_rdy | xls_float_ips__result_valid_inv;
  assign xls_float_ips__result_load_en = p0_all_active_inputs_valid & xls_float_ips__result_valid_load_en;
  assign nor_1037 = ~(and_1006 | and_1007 | (~(and_1006 | and_1007 | ~result) | nor_1012 & (eq_1002 & eq_exp & a_fraction__5 == b_fraction__2 | and_1009)));
  assign p0_stage_done = p0_all_active_inputs_valid & xls_float_ips__result_load_en;
  assign __xls_float_ips__result_buf = and_1006 | and_1007 | nor_1037;
  always @ (posedge clk) begin
    if (rst) begin
      __xls_float_ips__result_reg <= 1'h0;
      __xls_float_ips__result_valid_reg <= 1'h0;
    end else begin
      __xls_float_ips__result_reg <= xls_float_ips__result_load_en ? __xls_float_ips__result_buf : __xls_float_ips__result_reg;
      __xls_float_ips__result_valid_reg <= xls_float_ips__result_valid_load_en ? p0_all_active_inputs_valid : __xls_float_ips__result_valid_reg;
    end
  end
  assign xls_float_ips__result = __xls_float_ips__result_reg;
  assign xls_float_ips__result_vld = __xls_float_ips__result_valid_reg;
  assign xls_float_ips__lhs_rdy = p0_stage_done;
  assign xls_float_ips__rhs_rdy = p0_stage_done;
endmodule
module __xls_float_ips__divf32_0_next(
  input wire clk,
  input wire rst,
  input wire [31:0] xls_float_ips__lhs,
  input wire xls_float_ips__lhs_vld,
  input wire [31:0] xls_float_ips__rhs,
  input wire xls_float_ips__rhs_vld,
  input wire xls_float_ips__result_rdy,
  output wire [31:0] xls_float_ips__result,
  output wire xls_float_ips__result_vld,
  output wire xls_float_ips__lhs_rdy,
  output wire xls_float_ips__rhs_rdy
);
  wire [31:0] __xls_float_ips__result_reg_init = {1'h0, 8'h00, 23'h00_0000};
  reg p0_bit_slice_3995;
  reg p0_bit_slice_3996;
  reg p0_bit_slice_3997;
  reg p0_bit_slice_3998;
  reg p0_bit_slice_3999;
  reg p0_bit_slice_4000;
  reg p0_bit_slice_4001;
  reg p0_bit_slice_4002;
  reg p0_bit_slice_4003;
  reg p0_bit_slice_4004;
  reg p0_bit_slice_4005;
  reg p0_bit_slice_4006;
  reg p0_bit_slice_4007;
  reg p0_bit_slice_4008;
  reg p0_bit_slice_4009;
  reg p0_bit_slice_4010;
  reg p0_bit_slice_4011;
  reg p0_bit_slice_4012;
  reg p0_bit_slice_4013;
  reg p0_bit_slice_4014;
  reg p0_bit_slice_4015;
  reg [7:0] p0_a_bexp;
  reg p0_bit_slice_4017;
  reg p0_bit_slice_4018;
  reg p0_a_sign;
  reg [22:0] p1_concat_4081;
  reg [22:0] p1_b_fraction;
  reg p1_bit_slice_3996;
  reg p1_bit_slice_3997;
  reg p1_bit_slice_3998;
  reg p1_bit_slice_3999;
  reg p1_bit_slice_4000;
  reg p1_bit_slice_4001;
  reg p1_bit_slice_4002;
  reg p1_bit_slice_4003;
  reg p1_bit_slice_4004;
  reg p1_bit_slice_4005;
  reg p1_bit_slice_4006;
  reg p1_bit_slice_4007;
  reg p1_bit_slice_4008;
  reg p1_bit_slice_4009;
  reg p1_bit_slice_4010;
  reg p1_bit_slice_4011;
  reg p1_bit_slice_4012;
  reg p1_bit_slice_4013;
  reg p1_bit_slice_4014;
  reg p1_bit_slice_4015;
  reg [7:0] p1_a_bexp;
  reg [7:0] p1_b_bexp;
  reg p1_bit_slice_4017;
  reg p1_bit_slice_4018;
  reg p1_result_sign;
  reg [22:0] p2_b_fraction;
  reg p2_uge_4144;
  reg [23:0] p2_b_fractionivisor__1;
  reg [22:0] p2_concat_4151;
  reg p2_uge_4152;
  reg p2_bit_slice_3997;
  reg p2_bit_slice_3998;
  reg p2_bit_slice_3999;
  reg p2_bit_slice_4000;
  reg p2_bit_slice_4001;
  reg p2_bit_slice_4002;
  reg p2_bit_slice_4003;
  reg p2_bit_slice_4004;
  reg p2_bit_slice_4005;
  reg p2_bit_slice_4006;
  reg p2_bit_slice_4007;
  reg p2_bit_slice_4008;
  reg p2_bit_slice_4009;
  reg p2_bit_slice_4010;
  reg p2_bit_slice_4011;
  reg p2_bit_slice_4012;
  reg p2_bit_slice_4013;
  reg p2_bit_slice_4014;
  reg p2_bit_slice_4015;
  reg p2_bit_slice_4017;
  reg [8:0] p2_signed_exp_s9;
  reg p2_bit_slice_4018;
  reg p2_result_sign;
  reg [22:0] p3_b_fraction;
  reg p3_uge_4144;
  reg [23:0] p3_b_fractionivisor__1;
  reg p3_uge_4152;
  reg [22:0] p3_concat_4222;
  reg p3_uge_4223;
  reg p3_bit_slice_3998;
  reg p3_bit_slice_3999;
  reg p3_bit_slice_4000;
  reg p3_bit_slice_4001;
  reg p3_bit_slice_4002;
  reg p3_bit_slice_4003;
  reg p3_bit_slice_4004;
  reg p3_bit_slice_4005;
  reg p3_bit_slice_4006;
  reg p3_bit_slice_4007;
  reg p3_bit_slice_4008;
  reg p3_bit_slice_4009;
  reg p3_bit_slice_4010;
  reg p3_bit_slice_4011;
  reg p3_bit_slice_4012;
  reg p3_bit_slice_4013;
  reg p3_bit_slice_4014;
  reg p3_bit_slice_4015;
  reg p3_bit_slice_4017;
  reg p3_bit_slice_4018;
  reg p3_flag_zero;
  reg p3_result_sign;
  reg [7:0] p3_result_exp;
  reg [22:0] p4_b_fraction;
  reg p4_uge_4144;
  reg [23:0] p4_b_fractionivisor__1;
  reg p4_uge_4152;
  reg p4_uge_4223;
  reg [22:0] p4_concat_4297;
  reg p4_uge_4298;
  reg p4_bit_slice_3999;
  reg p4_bit_slice_4000;
  reg p4_bit_slice_4001;
  reg p4_bit_slice_4002;
  reg p4_bit_slice_4003;
  reg p4_bit_slice_4004;
  reg p4_bit_slice_4005;
  reg p4_bit_slice_4006;
  reg p4_bit_slice_4007;
  reg p4_bit_slice_4008;
  reg p4_bit_slice_4009;
  reg p4_bit_slice_4010;
  reg p4_bit_slice_4011;
  reg p4_bit_slice_4012;
  reg p4_bit_slice_4013;
  reg p4_bit_slice_4014;
  reg p4_bit_slice_4015;
  reg p4_bit_slice_4017;
  reg p4_bit_slice_4018;
  reg p4_flag_zero;
  reg p4_result_sign;
  reg [7:0] p4_result_exp;
  reg [22:0] p5_b_fraction;
  reg p5_uge_4144;
  reg [23:0] p5_b_fractionivisor__1;
  reg p5_uge_4152;
  reg p5_uge_4223;
  reg p5_uge_4298;
  reg [22:0] p5_concat_4363;
  reg p5_uge_4364;
  reg p5_bit_slice_4000;
  reg p5_bit_slice_4001;
  reg p5_bit_slice_4002;
  reg p5_bit_slice_4003;
  reg p5_bit_slice_4004;
  reg p5_bit_slice_4005;
  reg p5_bit_slice_4006;
  reg p5_bit_slice_4007;
  reg p5_bit_slice_4008;
  reg p5_bit_slice_4009;
  reg p5_bit_slice_4010;
  reg p5_bit_slice_4011;
  reg p5_bit_slice_4012;
  reg p5_bit_slice_4013;
  reg p5_bit_slice_4014;
  reg p5_bit_slice_4015;
  reg p5_bit_slice_4017;
  reg p5_bit_slice_4018;
  reg p5_flag_zero;
  reg p5_result_sign;
  reg [7:0] p5_result_exp;
  reg [22:0] p6_b_fraction;
  reg p6_uge_4144;
  reg [23:0] p6_b_fractionivisor__1;
  reg p6_uge_4152;
  reg p6_uge_4223;
  reg p6_uge_4298;
  reg p6_uge_4364;
  reg [22:0] p6_concat_4429;
  reg p6_uge_4430;
  reg p6_bit_slice_4001;
  reg p6_bit_slice_4002;
  reg p6_bit_slice_4003;
  reg p6_bit_slice_4004;
  reg p6_bit_slice_4005;
  reg p6_bit_slice_4006;
  reg p6_bit_slice_4007;
  reg p6_bit_slice_4008;
  reg p6_bit_slice_4009;
  reg p6_bit_slice_4010;
  reg p6_bit_slice_4011;
  reg p6_bit_slice_4012;
  reg p6_bit_slice_4013;
  reg p6_bit_slice_4014;
  reg p6_bit_slice_4015;
  reg p6_bit_slice_4017;
  reg p6_bit_slice_4018;
  reg p6_flag_zero;
  reg p6_result_sign;
  reg [7:0] p6_result_exp;
  reg [22:0] p7_b_fraction;
  reg p7_uge_4144;
  reg [23:0] p7_b_fractionivisor__1;
  reg p7_uge_4152;
  reg p7_uge_4223;
  reg p7_uge_4298;
  reg p7_uge_4364;
  reg p7_uge_4430;
  reg [22:0] p7_concat_4495;
  reg p7_uge_4496;
  reg p7_bit_slice_4002;
  reg p7_bit_slice_4003;
  reg p7_bit_slice_4004;
  reg p7_bit_slice_4005;
  reg p7_bit_slice_4006;
  reg p7_bit_slice_4007;
  reg p7_bit_slice_4008;
  reg p7_bit_slice_4009;
  reg p7_bit_slice_4010;
  reg p7_bit_slice_4011;
  reg p7_bit_slice_4012;
  reg p7_bit_slice_4013;
  reg p7_bit_slice_4014;
  reg p7_bit_slice_4015;
  reg p7_bit_slice_4017;
  reg p7_bit_slice_4018;
  reg p7_flag_zero;
  reg p7_result_sign;
  reg [7:0] p7_result_exp;
  reg [22:0] p8_b_fraction;
  reg p8_uge_4144;
  reg [23:0] p8_b_fractionivisor__1;
  reg p8_uge_4152;
  reg p8_uge_4223;
  reg p8_uge_4298;
  reg p8_uge_4364;
  reg p8_uge_4430;
  reg p8_uge_4496;
  reg [22:0] p8_concat_4561;
  reg p8_uge_4562;
  reg p8_bit_slice_4003;
  reg p8_bit_slice_4004;
  reg p8_bit_slice_4005;
  reg p8_bit_slice_4006;
  reg p8_bit_slice_4007;
  reg p8_bit_slice_4008;
  reg p8_bit_slice_4009;
  reg p8_bit_slice_4010;
  reg p8_bit_slice_4011;
  reg p8_bit_slice_4012;
  reg p8_bit_slice_4013;
  reg p8_bit_slice_4014;
  reg p8_bit_slice_4015;
  reg p8_bit_slice_4017;
  reg p8_bit_slice_4018;
  reg p8_flag_zero;
  reg p8_result_sign;
  reg [7:0] p8_result_exp;
  reg [22:0] p9_b_fraction;
  reg p9_uge_4144;
  reg [23:0] p9_b_fractionivisor__1;
  reg p9_uge_4152;
  reg p9_uge_4223;
  reg p9_uge_4298;
  reg p9_uge_4364;
  reg p9_uge_4430;
  reg p9_uge_4496;
  reg p9_uge_4562;
  reg [22:0] p9_concat_4627;
  reg p9_uge_4628;
  reg p9_bit_slice_4004;
  reg p9_bit_slice_4005;
  reg p9_bit_slice_4006;
  reg p9_bit_slice_4007;
  reg p9_bit_slice_4008;
  reg p9_bit_slice_4009;
  reg p9_bit_slice_4010;
  reg p9_bit_slice_4011;
  reg p9_bit_slice_4012;
  reg p9_bit_slice_4013;
  reg p9_bit_slice_4014;
  reg p9_bit_slice_4015;
  reg p9_bit_slice_4017;
  reg p9_bit_slice_4018;
  reg p9_flag_zero;
  reg p9_result_sign;
  reg [7:0] p9_result_exp;
  reg [22:0] p10_b_fraction;
  reg p10_uge_4144;
  reg [23:0] p10_b_fractionivisor__1;
  reg p10_uge_4152;
  reg p10_uge_4223;
  reg p10_uge_4298;
  reg p10_uge_4364;
  reg p10_uge_4430;
  reg p10_uge_4496;
  reg p10_uge_4562;
  reg p10_uge_4628;
  reg [22:0] p10_concat_4693;
  reg p10_uge_4694;
  reg p10_bit_slice_4005;
  reg p10_bit_slice_4006;
  reg p10_bit_slice_4007;
  reg p10_bit_slice_4008;
  reg p10_bit_slice_4009;
  reg p10_bit_slice_4010;
  reg p10_bit_slice_4011;
  reg p10_bit_slice_4012;
  reg p10_bit_slice_4013;
  reg p10_bit_slice_4014;
  reg p10_bit_slice_4015;
  reg p10_bit_slice_4017;
  reg p10_bit_slice_4018;
  reg p10_flag_zero;
  reg p10_result_sign;
  reg [7:0] p10_result_exp;
  reg [22:0] p11_b_fraction;
  reg p11_uge_4144;
  reg [23:0] p11_b_fractionivisor__1;
  reg p11_uge_4152;
  reg p11_uge_4223;
  reg p11_uge_4298;
  reg p11_uge_4364;
  reg p11_uge_4430;
  reg p11_uge_4496;
  reg p11_uge_4562;
  reg p11_uge_4628;
  reg p11_uge_4694;
  reg [22:0] p11_concat_4759;
  reg p11_uge_4760;
  reg p11_bit_slice_4006;
  reg p11_bit_slice_4007;
  reg p11_bit_slice_4008;
  reg p11_bit_slice_4009;
  reg p11_bit_slice_4010;
  reg p11_bit_slice_4011;
  reg p11_bit_slice_4012;
  reg p11_bit_slice_4013;
  reg p11_bit_slice_4014;
  reg p11_bit_slice_4015;
  reg p11_bit_slice_4017;
  reg p11_bit_slice_4018;
  reg p11_flag_zero;
  reg p11_result_sign;
  reg [7:0] p11_result_exp;
  reg [22:0] p12_b_fraction;
  reg p12_uge_4144;
  reg [23:0] p12_b_fractionivisor__1;
  reg p12_uge_4152;
  reg p12_uge_4223;
  reg p12_uge_4298;
  reg p12_uge_4364;
  reg p12_uge_4430;
  reg p12_uge_4496;
  reg p12_uge_4562;
  reg p12_uge_4628;
  reg p12_uge_4694;
  reg p12_uge_4760;
  reg [22:0] p12_concat_4825;
  reg p12_uge_4826;
  reg p12_bit_slice_4007;
  reg p12_bit_slice_4008;
  reg p12_bit_slice_4009;
  reg p12_bit_slice_4010;
  reg p12_bit_slice_4011;
  reg p12_bit_slice_4012;
  reg p12_bit_slice_4013;
  reg p12_bit_slice_4014;
  reg p12_bit_slice_4015;
  reg p12_bit_slice_4017;
  reg p12_bit_slice_4018;
  reg p12_flag_zero;
  reg p12_result_sign;
  reg [7:0] p12_result_exp;
  reg [22:0] p13_b_fraction;
  reg p13_uge_4144;
  reg [23:0] p13_b_fractionivisor__1;
  reg p13_uge_4152;
  reg p13_uge_4223;
  reg p13_uge_4298;
  reg p13_uge_4364;
  reg p13_uge_4430;
  reg p13_uge_4496;
  reg p13_uge_4562;
  reg p13_uge_4628;
  reg p13_uge_4694;
  reg p13_uge_4760;
  reg p13_uge_4826;
  reg [22:0] p13_concat_4891;
  reg p13_uge_4892;
  reg p13_bit_slice_4008;
  reg p13_bit_slice_4009;
  reg p13_bit_slice_4010;
  reg p13_bit_slice_4011;
  reg p13_bit_slice_4012;
  reg p13_bit_slice_4013;
  reg p13_bit_slice_4014;
  reg p13_bit_slice_4015;
  reg p13_bit_slice_4017;
  reg p13_bit_slice_4018;
  reg p13_flag_zero;
  reg p13_result_sign;
  reg [7:0] p13_result_exp;
  reg [22:0] p14_b_fraction;
  reg p14_uge_4144;
  reg [23:0] p14_b_fractionivisor__1;
  reg p14_uge_4152;
  reg p14_uge_4223;
  reg p14_uge_4298;
  reg p14_uge_4364;
  reg p14_uge_4430;
  reg p14_uge_4496;
  reg p14_uge_4562;
  reg p14_uge_4628;
  reg p14_uge_4694;
  reg p14_uge_4760;
  reg p14_uge_4826;
  reg p14_uge_4892;
  reg [22:0] p14_concat_4957;
  reg p14_uge_4958;
  reg p14_bit_slice_4009;
  reg p14_bit_slice_4010;
  reg p14_bit_slice_4011;
  reg p14_bit_slice_4012;
  reg p14_bit_slice_4013;
  reg p14_bit_slice_4014;
  reg p14_bit_slice_4015;
  reg p14_bit_slice_4017;
  reg p14_bit_slice_4018;
  reg p14_flag_zero;
  reg p14_result_sign;
  reg [7:0] p14_result_exp;
  reg [22:0] p15_b_fraction;
  reg p15_uge_4144;
  reg [23:0] p15_b_fractionivisor__1;
  reg p15_uge_4152;
  reg p15_uge_4223;
  reg p15_uge_4298;
  reg p15_uge_4364;
  reg p15_uge_4430;
  reg p15_uge_4496;
  reg p15_uge_4562;
  reg p15_uge_4628;
  reg p15_uge_4694;
  reg p15_uge_4760;
  reg p15_uge_4826;
  reg p15_uge_4892;
  reg p15_uge_4958;
  reg [22:0] p15_concat_5023;
  reg p15_uge_5024;
  reg p15_bit_slice_4010;
  reg p15_bit_slice_4011;
  reg p15_bit_slice_4012;
  reg p15_bit_slice_4013;
  reg p15_bit_slice_4014;
  reg p15_bit_slice_4015;
  reg p15_bit_slice_4017;
  reg p15_bit_slice_4018;
  reg p15_flag_zero;
  reg p15_result_sign;
  reg [7:0] p15_result_exp;
  reg [22:0] p16_b_fraction;
  reg p16_uge_4144;
  reg [23:0] p16_b_fractionivisor__1;
  reg p16_uge_4152;
  reg p16_uge_4223;
  reg p16_uge_4298;
  reg p16_uge_4364;
  reg p16_uge_4430;
  reg p16_uge_4496;
  reg p16_uge_4562;
  reg p16_uge_4628;
  reg p16_uge_4694;
  reg p16_uge_4760;
  reg p16_uge_4826;
  reg p16_uge_4892;
  reg p16_uge_4958;
  reg p16_uge_5024;
  reg [22:0] p16_concat_5089;
  reg p16_uge_5090;
  reg p16_bit_slice_4011;
  reg p16_bit_slice_4012;
  reg p16_bit_slice_4013;
  reg p16_bit_slice_4014;
  reg p16_bit_slice_4015;
  reg p16_bit_slice_4017;
  reg p16_bit_slice_4018;
  reg p16_flag_zero;
  reg p16_result_sign;
  reg [7:0] p16_result_exp;
  reg [22:0] p17_b_fraction;
  reg p17_uge_4144;
  reg [23:0] p17_b_fractionivisor__1;
  reg p17_uge_4152;
  reg p17_uge_4223;
  reg p17_uge_4298;
  reg p17_uge_4364;
  reg p17_uge_4430;
  reg p17_uge_4496;
  reg p17_uge_4562;
  reg p17_uge_4628;
  reg p17_uge_4694;
  reg p17_uge_4760;
  reg p17_uge_4826;
  reg p17_uge_4892;
  reg p17_uge_4958;
  reg p17_uge_5024;
  reg p17_uge_5090;
  reg [22:0] p17_concat_5155;
  reg p17_uge_5156;
  reg p17_bit_slice_4012;
  reg p17_bit_slice_4013;
  reg p17_bit_slice_4014;
  reg p17_bit_slice_4015;
  reg p17_bit_slice_4017;
  reg p17_bit_slice_4018;
  reg p17_flag_zero;
  reg p17_result_sign;
  reg [7:0] p17_result_exp;
  reg [22:0] p18_b_fraction;
  reg p18_uge_4144;
  reg [23:0] p18_b_fractionivisor__1;
  reg p18_uge_4152;
  reg p18_uge_4223;
  reg p18_uge_4298;
  reg p18_uge_4364;
  reg p18_uge_4430;
  reg p18_uge_4496;
  reg p18_uge_4562;
  reg p18_uge_4628;
  reg p18_uge_4694;
  reg p18_uge_4760;
  reg p18_uge_4826;
  reg p18_uge_4892;
  reg p18_uge_4958;
  reg p18_uge_5024;
  reg p18_uge_5090;
  reg p18_uge_5156;
  reg [22:0] p18_concat_5221;
  reg p18_uge_5222;
  reg p18_bit_slice_4013;
  reg p18_bit_slice_4014;
  reg p18_bit_slice_4015;
  reg p18_bit_slice_4017;
  reg p18_bit_slice_4018;
  reg p18_flag_zero;
  reg p18_result_sign;
  reg [7:0] p18_result_exp;
  reg [22:0] p19_b_fraction;
  reg p19_uge_4144;
  reg [23:0] p19_b_fractionivisor__1;
  reg p19_uge_4152;
  reg p19_uge_4223;
  reg p19_uge_4298;
  reg p19_uge_4364;
  reg p19_uge_4430;
  reg p19_uge_4496;
  reg p19_uge_4562;
  reg p19_uge_4628;
  reg p19_uge_4694;
  reg p19_uge_4760;
  reg p19_uge_4826;
  reg p19_uge_4892;
  reg p19_uge_4958;
  reg p19_uge_5024;
  reg p19_uge_5090;
  reg p19_uge_5156;
  reg p19_uge_5222;
  reg [22:0] p19_concat_5287;
  reg p19_uge_5288;
  reg p19_bit_slice_4014;
  reg p19_bit_slice_4015;
  reg p19_bit_slice_4017;
  reg p19_bit_slice_4018;
  reg p19_flag_zero;
  reg p19_result_sign;
  reg [7:0] p19_result_exp;
  reg [22:0] p20_b_fraction;
  reg p20_uge_4144;
  reg [23:0] p20_b_fractionivisor__1;
  reg p20_uge_4152;
  reg p20_uge_4223;
  reg p20_uge_4298;
  reg p20_uge_4364;
  reg p20_uge_4430;
  reg p20_uge_4496;
  reg p20_uge_4562;
  reg p20_uge_4628;
  reg p20_uge_4694;
  reg p20_uge_4760;
  reg p20_uge_4826;
  reg p20_uge_4892;
  reg p20_uge_4958;
  reg p20_uge_5024;
  reg p20_uge_5090;
  reg p20_uge_5156;
  reg p20_uge_5222;
  reg p20_uge_5288;
  reg [22:0] p20_concat_5353;
  reg p20_uge_5354;
  reg p20_bit_slice_4015;
  reg p20_bit_slice_4017;
  reg p20_bit_slice_4018;
  reg p20_flag_zero;
  reg p20_result_sign;
  reg [7:0] p20_result_exp;
  reg [22:0] p21_b_fraction;
  reg p21_uge_4144;
  reg [23:0] p21_b_fractionivisor__1;
  reg p21_uge_4152;
  reg p21_uge_4223;
  reg p21_uge_4298;
  reg p21_uge_4364;
  reg p21_uge_4430;
  reg p21_uge_4496;
  reg p21_uge_4562;
  reg p21_uge_4628;
  reg p21_uge_4694;
  reg p21_uge_4760;
  reg p21_uge_4826;
  reg p21_uge_4892;
  reg p21_uge_4958;
  reg p21_uge_5024;
  reg p21_uge_5090;
  reg p21_uge_5156;
  reg p21_uge_5222;
  reg p21_uge_5288;
  reg p21_uge_5354;
  reg [22:0] p21_concat_5419;
  reg p21_uge_5420;
  reg p21_bit_slice_4017;
  reg p21_bit_slice_4018;
  reg p21_flag_zero;
  reg p21_result_sign;
  reg [7:0] p21_result_exp;
  reg [22:0] p22_b_fraction;
  reg p22_uge_4144;
  reg [23:0] p22_b_fractionivisor__1;
  reg p22_uge_4152;
  reg p22_uge_4223;
  reg p22_uge_4298;
  reg p22_uge_4364;
  reg p22_uge_4430;
  reg p22_uge_4496;
  reg p22_uge_4562;
  reg p22_uge_4628;
  reg p22_uge_4694;
  reg p22_uge_4760;
  reg p22_uge_4826;
  reg p22_uge_4892;
  reg p22_uge_4958;
  reg p22_uge_5024;
  reg p22_uge_5090;
  reg p22_uge_5156;
  reg p22_uge_5222;
  reg p22_uge_5288;
  reg p22_uge_5354;
  reg p22_uge_5420;
  reg [22:0] p22_concat_5485;
  reg p22_uge_5486;
  reg p22_bit_slice_4018;
  reg p22_flag_zero;
  reg p22_result_sign;
  reg [7:0] p22_result_exp;
  reg p23_uge_4144;
  reg p23_uge_4152;
  reg p23_uge_4223;
  reg p23_uge_4298;
  reg p23_uge_4364;
  reg p23_uge_4430;
  reg p23_uge_4496;
  reg p23_uge_4562;
  reg p23_uge_4628;
  reg p23_uge_4694;
  reg p23_uge_4760;
  reg p23_uge_4826;
  reg p23_uge_4892;
  reg p23_uge_4958;
  reg p23_uge_5024;
  reg p23_uge_5090;
  reg p23_uge_5156;
  reg p23_uge_5222;
  reg p23_uge_5288;
  reg p23_uge_5354;
  reg p23_uge_5420;
  reg p23_uge_5486;
  reg p23_flag_zero;
  reg p23_q__23_squeezed_portion_0_width_1;
  reg p23_result_sign;
  reg [7:0] p23_result_exp;
  reg p0_valid;
  reg p1_valid;
  reg p2_valid;
  reg p3_valid;
  reg p4_valid;
  reg p5_valid;
  reg p6_valid;
  reg p7_valid;
  reg p8_valid;
  reg p9_valid;
  reg p10_valid;
  reg p11_valid;
  reg p12_valid;
  reg p13_valid;
  reg p14_valid;
  reg p15_valid;
  reg p16_valid;
  reg p17_valid;
  reg p18_valid;
  reg p19_valid;
  reg p20_valid;
  reg p21_valid;
  reg p22_valid;
  reg p23_valid;
  reg p24_valid;
  reg p25_valid;
  reg p26_valid;
  reg p27_valid;
  reg p28_valid;
  reg [31:0] __xls_float_ips__result_reg;
  reg __xls_float_ips__result_valid_reg;
  wire xls_float_ips__result_valid_inv;
  wire xls_float_ips__result_valid_load_en;
  wire xls_float_ips__result_load_en;
  wire p24_stage_done;
  wire p24_not_valid;
  wire p23_enable;
  wire p23_data_enable;
  wire p23_not_valid;
  wire p22_enable;
  wire p22_data_enable;
  wire p22_not_valid;
  wire p21_enable;
  wire p21_data_enable;
  wire p21_not_valid;
  wire p20_enable;
  wire p20_data_enable;
  wire p20_not_valid;
  wire p19_enable;
  wire p19_data_enable;
  wire p19_not_valid;
  wire p18_enable;
  wire p18_data_enable;
  wire p18_not_valid;
  wire p17_enable;
  wire p17_data_enable;
  wire p17_not_valid;
  wire p16_enable;
  wire p16_data_enable;
  wire p16_not_valid;
  wire p15_enable;
  wire p15_data_enable;
  wire p15_not_valid;
  wire p14_enable;
  wire p14_data_enable;
  wire p14_not_valid;
  wire p13_enable;
  wire p13_data_enable;
  wire p13_not_valid;
  wire p12_enable;
  wire p12_data_enable;
  wire p12_not_valid;
  wire p11_enable;
  wire p11_data_enable;
  wire p11_not_valid;
  wire p10_enable;
  wire p10_data_enable;
  wire p10_not_valid;
  wire p9_enable;
  wire p9_data_enable;
  wire p9_not_valid;
  wire p8_enable;
  wire p8_data_enable;
  wire p8_not_valid;
  wire p7_enable;
  wire p7_data_enable;
  wire p7_not_valid;
  wire p6_enable;
  wire p6_data_enable;
  wire p6_not_valid;
  wire p5_enable;
  wire p5_data_enable;
  wire p5_not_valid;
  wire p4_enable;
  wire p4_data_enable;
  wire p4_not_valid;
  wire p3_enable;
  wire p3_data_enable;
  wire p3_not_valid;
  wire p2_enable;
  wire p2_data_enable;
  wire p2_not_valid;
  wire [22:0] sub_5547;
  wire [22:0] sub_5481;
  wire [22:0] sub_5415;
  wire [22:0] sub_5349;
  wire [22:0] sub_5283;
  wire [22:0] sub_5217;
  wire [22:0] sub_5151;
  wire [22:0] sub_5085;
  wire [22:0] sub_5019;
  wire [22:0] sub_4953;
  wire [22:0] sub_4887;
  wire [22:0] sub_4821;
  wire [22:0] sub_4755;
  wire [22:0] sub_4689;
  wire [22:0] sub_4623;
  wire [22:0] sub_4557;
  wire [22:0] sub_4491;
  wire [22:0] sub_4425;
  wire [22:0] sub_4359;
  wire [22:0] sub_4293;
  wire [22:0] sub_4218;
  wire flag_zero;
  wire uge_4144;
  wire [22:0] sub_4145;
  wire p1_enable;
  wire p1_stage_done;
  wire [22:0] r__44;
  wire [22:0] r__42;
  wire [22:0] r__40;
  wire [22:0] r__38;
  wire [22:0] r__36;
  wire [22:0] r__34;
  wire [22:0] r__32;
  wire [22:0] r__30;
  wire [22:0] r__28;
  wire [22:0] r__26;
  wire [22:0] r__24;
  wire [22:0] r__22;
  wire [22:0] r__20;
  wire [22:0] r__18;
  wire [22:0] r__16;
  wire [22:0] r__14;
  wire [22:0] r__12;
  wire [22:0] r__10;
  wire [22:0] r__8;
  wire [22:0] r__6;
  wire [22:0] r__4;
  wire flag_inf;
  wire [22:0] r__2;
  wire p1_data_enable;
  wire p1_not_valid;
  wire [22:0] q__23;
  wire [23:0] r__45;
  wire [23:0] r__43;
  wire [23:0] r__41;
  wire [23:0] r__39;
  wire [23:0] r__37;
  wire [23:0] r__35;
  wire [23:0] r__33;
  wire [23:0] r__31;
  wire [23:0] r__29;
  wire [23:0] r__27;
  wire [23:0] r__25;
  wire [23:0] r__23;
  wire [23:0] r__21;
  wire [23:0] r__19;
  wire [23:0] r__17;
  wire [23:0] r__15;
  wire [23:0] r__13;
  wire [23:0] r__11;
  wire [23:0] r__9;
  wire [23:0] r__7;
  wire [23:0] r__5;
  wire [23:0] r__3;
  wire [23:0] b_fractionivisor__1;
  wire [8:0] sub_4157;
  wire b_sign;
  wire [22:0] a_fraction;
  wire p0_enable;
  wire [22:0] result_fraction;
  wire p28_enable;
  wire p27_enable;
  wire p26_enable;
  wire p25_enable;
  wire p24_enable;
  wire q__23_squeezed_portion_0_width_1;
  wire [22:0] concat_5485;
  wire uge_5486;
  wire [22:0] concat_5419;
  wire uge_5420;
  wire [22:0] concat_5353;
  wire uge_5354;
  wire [22:0] concat_5287;
  wire uge_5288;
  wire [22:0] concat_5221;
  wire uge_5222;
  wire [22:0] concat_5155;
  wire uge_5156;
  wire [22:0] concat_5089;
  wire uge_5090;
  wire [22:0] concat_5023;
  wire uge_5024;
  wire [22:0] concat_4957;
  wire uge_4958;
  wire [22:0] concat_4891;
  wire uge_4892;
  wire [22:0] concat_4825;
  wire uge_4826;
  wire [22:0] concat_4759;
  wire uge_4760;
  wire [22:0] concat_4693;
  wire uge_4694;
  wire [22:0] concat_4627;
  wire uge_4628;
  wire [22:0] concat_4561;
  wire uge_4562;
  wire [22:0] concat_4495;
  wire uge_4496;
  wire [22:0] concat_4429;
  wire uge_4430;
  wire [22:0] concat_4363;
  wire uge_4364;
  wire [22:0] concat_4297;
  wire uge_4298;
  wire [22:0] concat_4222;
  wire uge_4223;
  wire [7:0] result_exp;
  wire [22:0] concat_4151;
  wire uge_4152;
  wire [8:0] signed_exp_s9;
  wire [22:0] concat_4081;
  wire [22:0] b_fraction;
  wire [7:0] b_bexp;
  wire result_sign;
  wire bit_slice_3995;
  wire p0_data_enable;
  wire bit_slice_3996;
  wire bit_slice_3997;
  wire bit_slice_3998;
  wire bit_slice_3999;
  wire bit_slice_4000;
  wire bit_slice_4001;
  wire bit_slice_4002;
  wire bit_slice_4003;
  wire bit_slice_4004;
  wire bit_slice_4005;
  wire bit_slice_4006;
  wire bit_slice_4007;
  wire bit_slice_4008;
  wire bit_slice_4009;
  wire bit_slice_4010;
  wire bit_slice_4011;
  wire bit_slice_4012;
  wire bit_slice_4013;
  wire bit_slice_4014;
  wire bit_slice_4015;
  wire [7:0] a_bexp;
  wire bit_slice_4017;
  wire bit_slice_4018;
  wire a_sign;
  wire [31:0] __xls_float_ips__result_buf;
  assign xls_float_ips__result_valid_inv = ~__xls_float_ips__result_valid_reg;
  assign xls_float_ips__result_valid_load_en = xls_float_ips__result_rdy | xls_float_ips__result_valid_inv;
  assign xls_float_ips__result_load_en = p23_valid & xls_float_ips__result_valid_load_en;
  assign p24_stage_done = p23_valid & xls_float_ips__result_load_en;
  assign p24_not_valid = ~p23_valid;
  assign p23_enable = p24_stage_done | p24_not_valid;
  assign p23_data_enable = p23_enable & p22_valid;
  assign p23_not_valid = ~p22_valid;
  assign p22_enable = p23_data_enable | p23_not_valid;
  assign p22_data_enable = p22_enable & p21_valid;
  assign p22_not_valid = ~p21_valid;
  assign p21_enable = p22_data_enable | p22_not_valid;
  assign p21_data_enable = p21_enable & p20_valid;
  assign p21_not_valid = ~p20_valid;
  assign p20_enable = p21_data_enable | p21_not_valid;
  assign p20_data_enable = p20_enable & p19_valid;
  assign p20_not_valid = ~p19_valid;
  assign p19_enable = p20_data_enable | p20_not_valid;
  assign p19_data_enable = p19_enable & p18_valid;
  assign p19_not_valid = ~p18_valid;
  assign p18_enable = p19_data_enable | p19_not_valid;
  assign p18_data_enable = p18_enable & p17_valid;
  assign p18_not_valid = ~p17_valid;
  assign p17_enable = p18_data_enable | p18_not_valid;
  assign p17_data_enable = p17_enable & p16_valid;
  assign p17_not_valid = ~p16_valid;
  assign p16_enable = p17_data_enable | p17_not_valid;
  assign p16_data_enable = p16_enable & p15_valid;
  assign p16_not_valid = ~p15_valid;
  assign p15_enable = p16_data_enable | p16_not_valid;
  assign p15_data_enable = p15_enable & p14_valid;
  assign p15_not_valid = ~p14_valid;
  assign p14_enable = p15_data_enable | p15_not_valid;
  assign p14_data_enable = p14_enable & p13_valid;
  assign p14_not_valid = ~p13_valid;
  assign p13_enable = p14_data_enable | p14_not_valid;
  assign p13_data_enable = p13_enable & p12_valid;
  assign p13_not_valid = ~p12_valid;
  assign p12_enable = p13_data_enable | p13_not_valid;
  assign p12_data_enable = p12_enable & p11_valid;
  assign p12_not_valid = ~p11_valid;
  assign p11_enable = p12_data_enable | p12_not_valid;
  assign p11_data_enable = p11_enable & p10_valid;
  assign p11_not_valid = ~p10_valid;
  assign p10_enable = p11_data_enable | p11_not_valid;
  assign p10_data_enable = p10_enable & p9_valid;
  assign p10_not_valid = ~p9_valid;
  assign p9_enable = p10_data_enable | p10_not_valid;
  assign p9_data_enable = p9_enable & p8_valid;
  assign p9_not_valid = ~p8_valid;
  assign p8_enable = p9_data_enable | p9_not_valid;
  assign p8_data_enable = p8_enable & p7_valid;
  assign p8_not_valid = ~p7_valid;
  assign p7_enable = p8_data_enable | p8_not_valid;
  assign p7_data_enable = p7_enable & p6_valid;
  assign p7_not_valid = ~p6_valid;
  assign p6_enable = p7_data_enable | p7_not_valid;
  assign p6_data_enable = p6_enable & p5_valid;
  assign p6_not_valid = ~p5_valid;
  assign p5_enable = p6_data_enable | p6_not_valid;
  assign p5_data_enable = p5_enable & p4_valid;
  assign p5_not_valid = ~p4_valid;
  assign p4_enable = p5_data_enable | p5_not_valid;
  assign p4_data_enable = p4_enable & p3_valid;
  assign p4_not_valid = ~p3_valid;
  assign p3_enable = p4_data_enable | p4_not_valid;
  assign p3_data_enable = p3_enable & p2_valid;
  assign p3_not_valid = ~p2_valid;
  assign p2_enable = p3_data_enable | p3_not_valid;
  assign p2_data_enable = p2_enable & p1_valid;
  assign p2_not_valid = ~p1_valid;
  assign sub_5547 = p22_concat_5485 - p22_b_fraction;
  assign sub_5481 = p21_concat_5419 - p21_b_fraction;
  assign sub_5415 = p20_concat_5353 - p20_b_fraction;
  assign sub_5349 = p19_concat_5287 - p19_b_fraction;
  assign sub_5283 = p18_concat_5221 - p18_b_fraction;
  assign sub_5217 = p17_concat_5155 - p17_b_fraction;
  assign sub_5151 = p16_concat_5089 - p16_b_fraction;
  assign sub_5085 = p15_concat_5023 - p15_b_fraction;
  assign sub_5019 = p14_concat_4957 - p14_b_fraction;
  assign sub_4953 = p13_concat_4891 - p13_b_fraction;
  assign sub_4887 = p12_concat_4825 - p12_b_fraction;
  assign sub_4821 = p11_concat_4759 - p11_b_fraction;
  assign sub_4755 = p10_concat_4693 - p10_b_fraction;
  assign sub_4689 = p9_concat_4627 - p9_b_fraction;
  assign sub_4623 = p8_concat_4561 - p8_b_fraction;
  assign sub_4557 = p7_concat_4495 - p7_b_fraction;
  assign sub_4491 = p6_concat_4429 - p6_b_fraction;
  assign sub_4425 = p5_concat_4363 - p5_b_fraction;
  assign sub_4359 = p4_concat_4297 - p4_b_fraction;
  assign sub_4293 = p3_concat_4222 - p3_b_fraction;
  assign sub_4218 = p2_concat_4151 - p2_b_fraction;
  assign flag_zero = p2_signed_exp_s9[8];
  assign uge_4144 = p1_concat_4081 >= p1_b_fraction;
  assign sub_4145 = p1_concat_4081 - p1_b_fraction;
  assign p1_enable = p2_data_enable | p2_not_valid;
  assign p1_stage_done = p0_valid & xls_float_ips__rhs_vld;
  assign r__44 = p22_uge_5486 ? sub_5547 : p22_concat_5485;
  assign r__42 = p21_uge_5420 ? sub_5481 : p21_concat_5419;
  assign r__40 = p20_uge_5354 ? sub_5415 : p20_concat_5353;
  assign r__38 = p19_uge_5288 ? sub_5349 : p19_concat_5287;
  assign r__36 = p18_uge_5222 ? sub_5283 : p18_concat_5221;
  assign r__34 = p17_uge_5156 ? sub_5217 : p17_concat_5155;
  assign r__32 = p16_uge_5090 ? sub_5151 : p16_concat_5089;
  assign r__30 = p15_uge_5024 ? sub_5085 : p15_concat_5023;
  assign r__28 = p14_uge_4958 ? sub_5019 : p14_concat_4957;
  assign r__26 = p13_uge_4892 ? sub_4953 : p13_concat_4891;
  assign r__24 = p12_uge_4826 ? sub_4887 : p12_concat_4825;
  assign r__22 = p11_uge_4760 ? sub_4821 : p11_concat_4759;
  assign r__20 = p10_uge_4694 ? sub_4755 : p10_concat_4693;
  assign r__18 = p9_uge_4628 ? sub_4689 : p9_concat_4627;
  assign r__16 = p8_uge_4562 ? sub_4623 : p8_concat_4561;
  assign r__14 = p7_uge_4496 ? sub_4557 : p7_concat_4495;
  assign r__12 = p6_uge_4430 ? sub_4491 : p6_concat_4429;
  assign r__10 = p5_uge_4364 ? sub_4425 : p5_concat_4363;
  assign r__8 = p4_uge_4298 ? sub_4359 : p4_concat_4297;
  assign r__6 = p3_uge_4223 ? sub_4293 : p3_concat_4222;
  assign r__4 = p2_uge_4152 ? sub_4218 : p2_concat_4151;
  assign flag_inf = $signed(p2_signed_exp_s9) > $signed(9'h0fe);
  assign r__2 = uge_4144 ? sub_4145 : p1_concat_4081;
  assign p1_data_enable = p1_enable & p1_stage_done;
  assign p1_not_valid = ~p0_valid;
  assign q__23 = {p23_uge_4144, p23_uge_4152, p23_uge_4223, p23_uge_4298, p23_uge_4364, p23_uge_4430, p23_uge_4496, p23_uge_4562, p23_uge_4628, p23_uge_4694, p23_uge_4760, p23_uge_4826, p23_uge_4892, p23_uge_4958, p23_uge_5024, p23_uge_5090, p23_uge_5156, p23_uge_5222, p23_uge_5288, p23_uge_5354, p23_uge_5420, p23_uge_5486, p23_q__23_squeezed_portion_0_width_1};
  assign r__45 = {r__44, p22_bit_slice_4018};
  assign r__43 = {r__42, p21_bit_slice_4017};
  assign r__41 = {r__40, p20_bit_slice_4015};
  assign r__39 = {r__38, p19_bit_slice_4014};
  assign r__37 = {r__36, p18_bit_slice_4013};
  assign r__35 = {r__34, p17_bit_slice_4012};
  assign r__33 = {r__32, p16_bit_slice_4011};
  assign r__31 = {r__30, p15_bit_slice_4010};
  assign r__29 = {r__28, p14_bit_slice_4009};
  assign r__27 = {r__26, p13_bit_slice_4008};
  assign r__25 = {r__24, p12_bit_slice_4007};
  assign r__23 = {r__22, p11_bit_slice_4006};
  assign r__21 = {r__20, p10_bit_slice_4005};
  assign r__19 = {r__18, p9_bit_slice_4004};
  assign r__17 = {r__16, p8_bit_slice_4003};
  assign r__15 = {r__14, p7_bit_slice_4002};
  assign r__13 = {r__12, p6_bit_slice_4001};
  assign r__11 = {r__10, p5_bit_slice_4000};
  assign r__9 = {r__8, p4_bit_slice_3999};
  assign r__7 = {r__6, p3_bit_slice_3998};
  assign r__5 = {r__4, p2_bit_slice_3997};
  assign r__3 = {r__2, p1_bit_slice_3996};
  assign b_fractionivisor__1 = {1'h0, p1_b_fraction};
  assign sub_4157 = {1'h0, p1_a_bexp} - {1'h0, p1_b_bexp};
  assign b_sign = xls_float_ips__rhs[31:31];
  assign a_fraction = xls_float_ips__lhs[22:0];
  assign p0_enable = p1_data_enable | p1_not_valid;
  assign result_fraction = p23_flag_zero ? 23'h00_0001 : q__23;
  assign p28_enable = 1'h1;
  assign p27_enable = 1'h1;
  assign p26_enable = 1'h1;
  assign p25_enable = 1'h1;
  assign p24_enable = 1'h1;
  assign q__23_squeezed_portion_0_width_1 = r__45 >= p22_b_fractionivisor__1;
  assign concat_5485 = {r__42[21:0], p21_bit_slice_4017};
  assign uge_5486 = r__43 >= p21_b_fractionivisor__1;
  assign concat_5419 = {r__40[21:0], p20_bit_slice_4015};
  assign uge_5420 = r__41 >= p20_b_fractionivisor__1;
  assign concat_5353 = {r__38[21:0], p19_bit_slice_4014};
  assign uge_5354 = r__39 >= p19_b_fractionivisor__1;
  assign concat_5287 = {r__36[21:0], p18_bit_slice_4013};
  assign uge_5288 = r__37 >= p18_b_fractionivisor__1;
  assign concat_5221 = {r__34[21:0], p17_bit_slice_4012};
  assign uge_5222 = r__35 >= p17_b_fractionivisor__1;
  assign concat_5155 = {r__32[21:0], p16_bit_slice_4011};
  assign uge_5156 = r__33 >= p16_b_fractionivisor__1;
  assign concat_5089 = {r__30[21:0], p15_bit_slice_4010};
  assign uge_5090 = r__31 >= p15_b_fractionivisor__1;
  assign concat_5023 = {r__28[21:0], p14_bit_slice_4009};
  assign uge_5024 = r__29 >= p14_b_fractionivisor__1;
  assign concat_4957 = {r__26[21:0], p13_bit_slice_4008};
  assign uge_4958 = r__27 >= p13_b_fractionivisor__1;
  assign concat_4891 = {r__24[21:0], p12_bit_slice_4007};
  assign uge_4892 = r__25 >= p12_b_fractionivisor__1;
  assign concat_4825 = {r__22[21:0], p11_bit_slice_4006};
  assign uge_4826 = r__23 >= p11_b_fractionivisor__1;
  assign concat_4759 = {r__20[21:0], p10_bit_slice_4005};
  assign uge_4760 = r__21 >= p10_b_fractionivisor__1;
  assign concat_4693 = {r__18[21:0], p9_bit_slice_4004};
  assign uge_4694 = r__19 >= p9_b_fractionivisor__1;
  assign concat_4627 = {r__16[21:0], p8_bit_slice_4003};
  assign uge_4628 = r__17 >= p8_b_fractionivisor__1;
  assign concat_4561 = {r__14[21:0], p7_bit_slice_4002};
  assign uge_4562 = r__15 >= p7_b_fractionivisor__1;
  assign concat_4495 = {r__12[21:0], p6_bit_slice_4001};
  assign uge_4496 = r__13 >= p6_b_fractionivisor__1;
  assign concat_4429 = {r__10[21:0], p5_bit_slice_4000};
  assign uge_4430 = r__11 >= p5_b_fractionivisor__1;
  assign concat_4363 = {r__8[21:0], p4_bit_slice_3999};
  assign uge_4364 = r__9 >= p4_b_fractionivisor__1;
  assign concat_4297 = {r__6[21:0], p3_bit_slice_3998};
  assign uge_4298 = r__7 >= p3_b_fractionivisor__1;
  assign concat_4222 = {r__4[21:0], p2_bit_slice_3997};
  assign uge_4223 = r__5 >= p2_b_fractionivisor__1;
  assign result_exp = (flag_inf ? 8'hff : p2_signed_exp_s9[7:0]) & {8{~flag_zero}};
  assign concat_4151 = {r__2[21:0], p1_bit_slice_3996};
  assign uge_4152 = r__3 >= b_fractionivisor__1;
  assign signed_exp_s9 = sub_4157 + 9'h07f;
  assign concat_4081 = {22'h00_0000, p0_bit_slice_3995};
  assign b_fraction = xls_float_ips__rhs[22:0];
  assign b_bexp = xls_float_ips__rhs[30:23];
  assign result_sign = p0_a_sign ^ b_sign;
  assign bit_slice_3995 = a_fraction[22];
  assign p0_data_enable = p0_enable & xls_float_ips__lhs_vld;
  assign bit_slice_3996 = a_fraction[21];
  assign bit_slice_3997 = a_fraction[20];
  assign bit_slice_3998 = a_fraction[19];
  assign bit_slice_3999 = a_fraction[18];
  assign bit_slice_4000 = a_fraction[17];
  assign bit_slice_4001 = a_fraction[16];
  assign bit_slice_4002 = a_fraction[15];
  assign bit_slice_4003 = a_fraction[14];
  assign bit_slice_4004 = a_fraction[13];
  assign bit_slice_4005 = a_fraction[12];
  assign bit_slice_4006 = a_fraction[11];
  assign bit_slice_4007 = a_fraction[10];
  assign bit_slice_4008 = a_fraction[9];
  assign bit_slice_4009 = a_fraction[8];
  assign bit_slice_4010 = a_fraction[7];
  assign bit_slice_4011 = a_fraction[6];
  assign bit_slice_4012 = a_fraction[5];
  assign bit_slice_4013 = a_fraction[4];
  assign bit_slice_4014 = a_fraction[3];
  assign bit_slice_4015 = a_fraction[2];
  assign a_bexp = xls_float_ips__lhs[30:23];
  assign bit_slice_4017 = a_fraction[1];
  assign bit_slice_4018 = a_fraction[0];
  assign a_sign = xls_float_ips__lhs[31:31];
  assign __xls_float_ips__result_buf = {p23_result_sign, p23_result_exp, result_fraction};
  always @ (posedge clk) begin
    if (rst) begin
      p0_bit_slice_3995 <= 1'h0;
      p0_bit_slice_3996 <= 1'h0;
      p0_bit_slice_3997 <= 1'h0;
      p0_bit_slice_3998 <= 1'h0;
      p0_bit_slice_3999 <= 1'h0;
      p0_bit_slice_4000 <= 1'h0;
      p0_bit_slice_4001 <= 1'h0;
      p0_bit_slice_4002 <= 1'h0;
      p0_bit_slice_4003 <= 1'h0;
      p0_bit_slice_4004 <= 1'h0;
      p0_bit_slice_4005 <= 1'h0;
      p0_bit_slice_4006 <= 1'h0;
      p0_bit_slice_4007 <= 1'h0;
      p0_bit_slice_4008 <= 1'h0;
      p0_bit_slice_4009 <= 1'h0;
      p0_bit_slice_4010 <= 1'h0;
      p0_bit_slice_4011 <= 1'h0;
      p0_bit_slice_4012 <= 1'h0;
      p0_bit_slice_4013 <= 1'h0;
      p0_bit_slice_4014 <= 1'h0;
      p0_bit_slice_4015 <= 1'h0;
      p0_a_bexp <= 8'h00;
      p0_bit_slice_4017 <= 1'h0;
      p0_bit_slice_4018 <= 1'h0;
      p0_a_sign <= 1'h0;
      p1_concat_4081 <= 23'h00_0000;
      p1_b_fraction <= 23'h00_0000;
      p1_bit_slice_3996 <= 1'h0;
      p1_bit_slice_3997 <= 1'h0;
      p1_bit_slice_3998 <= 1'h0;
      p1_bit_slice_3999 <= 1'h0;
      p1_bit_slice_4000 <= 1'h0;
      p1_bit_slice_4001 <= 1'h0;
      p1_bit_slice_4002 <= 1'h0;
      p1_bit_slice_4003 <= 1'h0;
      p1_bit_slice_4004 <= 1'h0;
      p1_bit_slice_4005 <= 1'h0;
      p1_bit_slice_4006 <= 1'h0;
      p1_bit_slice_4007 <= 1'h0;
      p1_bit_slice_4008 <= 1'h0;
      p1_bit_slice_4009 <= 1'h0;
      p1_bit_slice_4010 <= 1'h0;
      p1_bit_slice_4011 <= 1'h0;
      p1_bit_slice_4012 <= 1'h0;
      p1_bit_slice_4013 <= 1'h0;
      p1_bit_slice_4014 <= 1'h0;
      p1_bit_slice_4015 <= 1'h0;
      p1_a_bexp <= 8'h00;
      p1_b_bexp <= 8'h00;
      p1_bit_slice_4017 <= 1'h0;
      p1_bit_slice_4018 <= 1'h0;
      p1_result_sign <= 1'h0;
      p2_b_fraction <= 23'h00_0000;
      p2_uge_4144 <= 1'h0;
      p2_b_fractionivisor__1 <= 24'h00_0000;
      p2_concat_4151 <= 23'h00_0000;
      p2_uge_4152 <= 1'h0;
      p2_bit_slice_3997 <= 1'h0;
      p2_bit_slice_3998 <= 1'h0;
      p2_bit_slice_3999 <= 1'h0;
      p2_bit_slice_4000 <= 1'h0;
      p2_bit_slice_4001 <= 1'h0;
      p2_bit_slice_4002 <= 1'h0;
      p2_bit_slice_4003 <= 1'h0;
      p2_bit_slice_4004 <= 1'h0;
      p2_bit_slice_4005 <= 1'h0;
      p2_bit_slice_4006 <= 1'h0;
      p2_bit_slice_4007 <= 1'h0;
      p2_bit_slice_4008 <= 1'h0;
      p2_bit_slice_4009 <= 1'h0;
      p2_bit_slice_4010 <= 1'h0;
      p2_bit_slice_4011 <= 1'h0;
      p2_bit_slice_4012 <= 1'h0;
      p2_bit_slice_4013 <= 1'h0;
      p2_bit_slice_4014 <= 1'h0;
      p2_bit_slice_4015 <= 1'h0;
      p2_bit_slice_4017 <= 1'h0;
      p2_signed_exp_s9 <= 9'h000;
      p2_bit_slice_4018 <= 1'h0;
      p2_result_sign <= 1'h0;
      p3_b_fraction <= 23'h00_0000;
      p3_uge_4144 <= 1'h0;
      p3_b_fractionivisor__1 <= 24'h00_0000;
      p3_uge_4152 <= 1'h0;
      p3_concat_4222 <= 23'h00_0000;
      p3_uge_4223 <= 1'h0;
      p3_bit_slice_3998 <= 1'h0;
      p3_bit_slice_3999 <= 1'h0;
      p3_bit_slice_4000 <= 1'h0;
      p3_bit_slice_4001 <= 1'h0;
      p3_bit_slice_4002 <= 1'h0;
      p3_bit_slice_4003 <= 1'h0;
      p3_bit_slice_4004 <= 1'h0;
      p3_bit_slice_4005 <= 1'h0;
      p3_bit_slice_4006 <= 1'h0;
      p3_bit_slice_4007 <= 1'h0;
      p3_bit_slice_4008 <= 1'h0;
      p3_bit_slice_4009 <= 1'h0;
      p3_bit_slice_4010 <= 1'h0;
      p3_bit_slice_4011 <= 1'h0;
      p3_bit_slice_4012 <= 1'h0;
      p3_bit_slice_4013 <= 1'h0;
      p3_bit_slice_4014 <= 1'h0;
      p3_bit_slice_4015 <= 1'h0;
      p3_bit_slice_4017 <= 1'h0;
      p3_bit_slice_4018 <= 1'h0;
      p3_flag_zero <= 1'h0;
      p3_result_sign <= 1'h0;
      p3_result_exp <= 8'h00;
      p4_b_fraction <= 23'h00_0000;
      p4_uge_4144 <= 1'h0;
      p4_b_fractionivisor__1 <= 24'h00_0000;
      p4_uge_4152 <= 1'h0;
      p4_uge_4223 <= 1'h0;
      p4_concat_4297 <= 23'h00_0000;
      p4_uge_4298 <= 1'h0;
      p4_bit_slice_3999 <= 1'h0;
      p4_bit_slice_4000 <= 1'h0;
      p4_bit_slice_4001 <= 1'h0;
      p4_bit_slice_4002 <= 1'h0;
      p4_bit_slice_4003 <= 1'h0;
      p4_bit_slice_4004 <= 1'h0;
      p4_bit_slice_4005 <= 1'h0;
      p4_bit_slice_4006 <= 1'h0;
      p4_bit_slice_4007 <= 1'h0;
      p4_bit_slice_4008 <= 1'h0;
      p4_bit_slice_4009 <= 1'h0;
      p4_bit_slice_4010 <= 1'h0;
      p4_bit_slice_4011 <= 1'h0;
      p4_bit_slice_4012 <= 1'h0;
      p4_bit_slice_4013 <= 1'h0;
      p4_bit_slice_4014 <= 1'h0;
      p4_bit_slice_4015 <= 1'h0;
      p4_bit_slice_4017 <= 1'h0;
      p4_bit_slice_4018 <= 1'h0;
      p4_flag_zero <= 1'h0;
      p4_result_sign <= 1'h0;
      p4_result_exp <= 8'h00;
      p5_b_fraction <= 23'h00_0000;
      p5_uge_4144 <= 1'h0;
      p5_b_fractionivisor__1 <= 24'h00_0000;
      p5_uge_4152 <= 1'h0;
      p5_uge_4223 <= 1'h0;
      p5_uge_4298 <= 1'h0;
      p5_concat_4363 <= 23'h00_0000;
      p5_uge_4364 <= 1'h0;
      p5_bit_slice_4000 <= 1'h0;
      p5_bit_slice_4001 <= 1'h0;
      p5_bit_slice_4002 <= 1'h0;
      p5_bit_slice_4003 <= 1'h0;
      p5_bit_slice_4004 <= 1'h0;
      p5_bit_slice_4005 <= 1'h0;
      p5_bit_slice_4006 <= 1'h0;
      p5_bit_slice_4007 <= 1'h0;
      p5_bit_slice_4008 <= 1'h0;
      p5_bit_slice_4009 <= 1'h0;
      p5_bit_slice_4010 <= 1'h0;
      p5_bit_slice_4011 <= 1'h0;
      p5_bit_slice_4012 <= 1'h0;
      p5_bit_slice_4013 <= 1'h0;
      p5_bit_slice_4014 <= 1'h0;
      p5_bit_slice_4015 <= 1'h0;
      p5_bit_slice_4017 <= 1'h0;
      p5_bit_slice_4018 <= 1'h0;
      p5_flag_zero <= 1'h0;
      p5_result_sign <= 1'h0;
      p5_result_exp <= 8'h00;
      p6_b_fraction <= 23'h00_0000;
      p6_uge_4144 <= 1'h0;
      p6_b_fractionivisor__1 <= 24'h00_0000;
      p6_uge_4152 <= 1'h0;
      p6_uge_4223 <= 1'h0;
      p6_uge_4298 <= 1'h0;
      p6_uge_4364 <= 1'h0;
      p6_concat_4429 <= 23'h00_0000;
      p6_uge_4430 <= 1'h0;
      p6_bit_slice_4001 <= 1'h0;
      p6_bit_slice_4002 <= 1'h0;
      p6_bit_slice_4003 <= 1'h0;
      p6_bit_slice_4004 <= 1'h0;
      p6_bit_slice_4005 <= 1'h0;
      p6_bit_slice_4006 <= 1'h0;
      p6_bit_slice_4007 <= 1'h0;
      p6_bit_slice_4008 <= 1'h0;
      p6_bit_slice_4009 <= 1'h0;
      p6_bit_slice_4010 <= 1'h0;
      p6_bit_slice_4011 <= 1'h0;
      p6_bit_slice_4012 <= 1'h0;
      p6_bit_slice_4013 <= 1'h0;
      p6_bit_slice_4014 <= 1'h0;
      p6_bit_slice_4015 <= 1'h0;
      p6_bit_slice_4017 <= 1'h0;
      p6_bit_slice_4018 <= 1'h0;
      p6_flag_zero <= 1'h0;
      p6_result_sign <= 1'h0;
      p6_result_exp <= 8'h00;
      p7_b_fraction <= 23'h00_0000;
      p7_uge_4144 <= 1'h0;
      p7_b_fractionivisor__1 <= 24'h00_0000;
      p7_uge_4152 <= 1'h0;
      p7_uge_4223 <= 1'h0;
      p7_uge_4298 <= 1'h0;
      p7_uge_4364 <= 1'h0;
      p7_uge_4430 <= 1'h0;
      p7_concat_4495 <= 23'h00_0000;
      p7_uge_4496 <= 1'h0;
      p7_bit_slice_4002 <= 1'h0;
      p7_bit_slice_4003 <= 1'h0;
      p7_bit_slice_4004 <= 1'h0;
      p7_bit_slice_4005 <= 1'h0;
      p7_bit_slice_4006 <= 1'h0;
      p7_bit_slice_4007 <= 1'h0;
      p7_bit_slice_4008 <= 1'h0;
      p7_bit_slice_4009 <= 1'h0;
      p7_bit_slice_4010 <= 1'h0;
      p7_bit_slice_4011 <= 1'h0;
      p7_bit_slice_4012 <= 1'h0;
      p7_bit_slice_4013 <= 1'h0;
      p7_bit_slice_4014 <= 1'h0;
      p7_bit_slice_4015 <= 1'h0;
      p7_bit_slice_4017 <= 1'h0;
      p7_bit_slice_4018 <= 1'h0;
      p7_flag_zero <= 1'h0;
      p7_result_sign <= 1'h0;
      p7_result_exp <= 8'h00;
      p8_b_fraction <= 23'h00_0000;
      p8_uge_4144 <= 1'h0;
      p8_b_fractionivisor__1 <= 24'h00_0000;
      p8_uge_4152 <= 1'h0;
      p8_uge_4223 <= 1'h0;
      p8_uge_4298 <= 1'h0;
      p8_uge_4364 <= 1'h0;
      p8_uge_4430 <= 1'h0;
      p8_uge_4496 <= 1'h0;
      p8_concat_4561 <= 23'h00_0000;
      p8_uge_4562 <= 1'h0;
      p8_bit_slice_4003 <= 1'h0;
      p8_bit_slice_4004 <= 1'h0;
      p8_bit_slice_4005 <= 1'h0;
      p8_bit_slice_4006 <= 1'h0;
      p8_bit_slice_4007 <= 1'h0;
      p8_bit_slice_4008 <= 1'h0;
      p8_bit_slice_4009 <= 1'h0;
      p8_bit_slice_4010 <= 1'h0;
      p8_bit_slice_4011 <= 1'h0;
      p8_bit_slice_4012 <= 1'h0;
      p8_bit_slice_4013 <= 1'h0;
      p8_bit_slice_4014 <= 1'h0;
      p8_bit_slice_4015 <= 1'h0;
      p8_bit_slice_4017 <= 1'h0;
      p8_bit_slice_4018 <= 1'h0;
      p8_flag_zero <= 1'h0;
      p8_result_sign <= 1'h0;
      p8_result_exp <= 8'h00;
      p9_b_fraction <= 23'h00_0000;
      p9_uge_4144 <= 1'h0;
      p9_b_fractionivisor__1 <= 24'h00_0000;
      p9_uge_4152 <= 1'h0;
      p9_uge_4223 <= 1'h0;
      p9_uge_4298 <= 1'h0;
      p9_uge_4364 <= 1'h0;
      p9_uge_4430 <= 1'h0;
      p9_uge_4496 <= 1'h0;
      p9_uge_4562 <= 1'h0;
      p9_concat_4627 <= 23'h00_0000;
      p9_uge_4628 <= 1'h0;
      p9_bit_slice_4004 <= 1'h0;
      p9_bit_slice_4005 <= 1'h0;
      p9_bit_slice_4006 <= 1'h0;
      p9_bit_slice_4007 <= 1'h0;
      p9_bit_slice_4008 <= 1'h0;
      p9_bit_slice_4009 <= 1'h0;
      p9_bit_slice_4010 <= 1'h0;
      p9_bit_slice_4011 <= 1'h0;
      p9_bit_slice_4012 <= 1'h0;
      p9_bit_slice_4013 <= 1'h0;
      p9_bit_slice_4014 <= 1'h0;
      p9_bit_slice_4015 <= 1'h0;
      p9_bit_slice_4017 <= 1'h0;
      p9_bit_slice_4018 <= 1'h0;
      p9_flag_zero <= 1'h0;
      p9_result_sign <= 1'h0;
      p9_result_exp <= 8'h00;
      p10_b_fraction <= 23'h00_0000;
      p10_uge_4144 <= 1'h0;
      p10_b_fractionivisor__1 <= 24'h00_0000;
      p10_uge_4152 <= 1'h0;
      p10_uge_4223 <= 1'h0;
      p10_uge_4298 <= 1'h0;
      p10_uge_4364 <= 1'h0;
      p10_uge_4430 <= 1'h0;
      p10_uge_4496 <= 1'h0;
      p10_uge_4562 <= 1'h0;
      p10_uge_4628 <= 1'h0;
      p10_concat_4693 <= 23'h00_0000;
      p10_uge_4694 <= 1'h0;
      p10_bit_slice_4005 <= 1'h0;
      p10_bit_slice_4006 <= 1'h0;
      p10_bit_slice_4007 <= 1'h0;
      p10_bit_slice_4008 <= 1'h0;
      p10_bit_slice_4009 <= 1'h0;
      p10_bit_slice_4010 <= 1'h0;
      p10_bit_slice_4011 <= 1'h0;
      p10_bit_slice_4012 <= 1'h0;
      p10_bit_slice_4013 <= 1'h0;
      p10_bit_slice_4014 <= 1'h0;
      p10_bit_slice_4015 <= 1'h0;
      p10_bit_slice_4017 <= 1'h0;
      p10_bit_slice_4018 <= 1'h0;
      p10_flag_zero <= 1'h0;
      p10_result_sign <= 1'h0;
      p10_result_exp <= 8'h00;
      p11_b_fraction <= 23'h00_0000;
      p11_uge_4144 <= 1'h0;
      p11_b_fractionivisor__1 <= 24'h00_0000;
      p11_uge_4152 <= 1'h0;
      p11_uge_4223 <= 1'h0;
      p11_uge_4298 <= 1'h0;
      p11_uge_4364 <= 1'h0;
      p11_uge_4430 <= 1'h0;
      p11_uge_4496 <= 1'h0;
      p11_uge_4562 <= 1'h0;
      p11_uge_4628 <= 1'h0;
      p11_uge_4694 <= 1'h0;
      p11_concat_4759 <= 23'h00_0000;
      p11_uge_4760 <= 1'h0;
      p11_bit_slice_4006 <= 1'h0;
      p11_bit_slice_4007 <= 1'h0;
      p11_bit_slice_4008 <= 1'h0;
      p11_bit_slice_4009 <= 1'h0;
      p11_bit_slice_4010 <= 1'h0;
      p11_bit_slice_4011 <= 1'h0;
      p11_bit_slice_4012 <= 1'h0;
      p11_bit_slice_4013 <= 1'h0;
      p11_bit_slice_4014 <= 1'h0;
      p11_bit_slice_4015 <= 1'h0;
      p11_bit_slice_4017 <= 1'h0;
      p11_bit_slice_4018 <= 1'h0;
      p11_flag_zero <= 1'h0;
      p11_result_sign <= 1'h0;
      p11_result_exp <= 8'h00;
      p12_b_fraction <= 23'h00_0000;
      p12_uge_4144 <= 1'h0;
      p12_b_fractionivisor__1 <= 24'h00_0000;
      p12_uge_4152 <= 1'h0;
      p12_uge_4223 <= 1'h0;
      p12_uge_4298 <= 1'h0;
      p12_uge_4364 <= 1'h0;
      p12_uge_4430 <= 1'h0;
      p12_uge_4496 <= 1'h0;
      p12_uge_4562 <= 1'h0;
      p12_uge_4628 <= 1'h0;
      p12_uge_4694 <= 1'h0;
      p12_uge_4760 <= 1'h0;
      p12_concat_4825 <= 23'h00_0000;
      p12_uge_4826 <= 1'h0;
      p12_bit_slice_4007 <= 1'h0;
      p12_bit_slice_4008 <= 1'h0;
      p12_bit_slice_4009 <= 1'h0;
      p12_bit_slice_4010 <= 1'h0;
      p12_bit_slice_4011 <= 1'h0;
      p12_bit_slice_4012 <= 1'h0;
      p12_bit_slice_4013 <= 1'h0;
      p12_bit_slice_4014 <= 1'h0;
      p12_bit_slice_4015 <= 1'h0;
      p12_bit_slice_4017 <= 1'h0;
      p12_bit_slice_4018 <= 1'h0;
      p12_flag_zero <= 1'h0;
      p12_result_sign <= 1'h0;
      p12_result_exp <= 8'h00;
      p13_b_fraction <= 23'h00_0000;
      p13_uge_4144 <= 1'h0;
      p13_b_fractionivisor__1 <= 24'h00_0000;
      p13_uge_4152 <= 1'h0;
      p13_uge_4223 <= 1'h0;
      p13_uge_4298 <= 1'h0;
      p13_uge_4364 <= 1'h0;
      p13_uge_4430 <= 1'h0;
      p13_uge_4496 <= 1'h0;
      p13_uge_4562 <= 1'h0;
      p13_uge_4628 <= 1'h0;
      p13_uge_4694 <= 1'h0;
      p13_uge_4760 <= 1'h0;
      p13_uge_4826 <= 1'h0;
      p13_concat_4891 <= 23'h00_0000;
      p13_uge_4892 <= 1'h0;
      p13_bit_slice_4008 <= 1'h0;
      p13_bit_slice_4009 <= 1'h0;
      p13_bit_slice_4010 <= 1'h0;
      p13_bit_slice_4011 <= 1'h0;
      p13_bit_slice_4012 <= 1'h0;
      p13_bit_slice_4013 <= 1'h0;
      p13_bit_slice_4014 <= 1'h0;
      p13_bit_slice_4015 <= 1'h0;
      p13_bit_slice_4017 <= 1'h0;
      p13_bit_slice_4018 <= 1'h0;
      p13_flag_zero <= 1'h0;
      p13_result_sign <= 1'h0;
      p13_result_exp <= 8'h00;
      p14_b_fraction <= 23'h00_0000;
      p14_uge_4144 <= 1'h0;
      p14_b_fractionivisor__1 <= 24'h00_0000;
      p14_uge_4152 <= 1'h0;
      p14_uge_4223 <= 1'h0;
      p14_uge_4298 <= 1'h0;
      p14_uge_4364 <= 1'h0;
      p14_uge_4430 <= 1'h0;
      p14_uge_4496 <= 1'h0;
      p14_uge_4562 <= 1'h0;
      p14_uge_4628 <= 1'h0;
      p14_uge_4694 <= 1'h0;
      p14_uge_4760 <= 1'h0;
      p14_uge_4826 <= 1'h0;
      p14_uge_4892 <= 1'h0;
      p14_concat_4957 <= 23'h00_0000;
      p14_uge_4958 <= 1'h0;
      p14_bit_slice_4009 <= 1'h0;
      p14_bit_slice_4010 <= 1'h0;
      p14_bit_slice_4011 <= 1'h0;
      p14_bit_slice_4012 <= 1'h0;
      p14_bit_slice_4013 <= 1'h0;
      p14_bit_slice_4014 <= 1'h0;
      p14_bit_slice_4015 <= 1'h0;
      p14_bit_slice_4017 <= 1'h0;
      p14_bit_slice_4018 <= 1'h0;
      p14_flag_zero <= 1'h0;
      p14_result_sign <= 1'h0;
      p14_result_exp <= 8'h00;
      p15_b_fraction <= 23'h00_0000;
      p15_uge_4144 <= 1'h0;
      p15_b_fractionivisor__1 <= 24'h00_0000;
      p15_uge_4152 <= 1'h0;
      p15_uge_4223 <= 1'h0;
      p15_uge_4298 <= 1'h0;
      p15_uge_4364 <= 1'h0;
      p15_uge_4430 <= 1'h0;
      p15_uge_4496 <= 1'h0;
      p15_uge_4562 <= 1'h0;
      p15_uge_4628 <= 1'h0;
      p15_uge_4694 <= 1'h0;
      p15_uge_4760 <= 1'h0;
      p15_uge_4826 <= 1'h0;
      p15_uge_4892 <= 1'h0;
      p15_uge_4958 <= 1'h0;
      p15_concat_5023 <= 23'h00_0000;
      p15_uge_5024 <= 1'h0;
      p15_bit_slice_4010 <= 1'h0;
      p15_bit_slice_4011 <= 1'h0;
      p15_bit_slice_4012 <= 1'h0;
      p15_bit_slice_4013 <= 1'h0;
      p15_bit_slice_4014 <= 1'h0;
      p15_bit_slice_4015 <= 1'h0;
      p15_bit_slice_4017 <= 1'h0;
      p15_bit_slice_4018 <= 1'h0;
      p15_flag_zero <= 1'h0;
      p15_result_sign <= 1'h0;
      p15_result_exp <= 8'h00;
      p16_b_fraction <= 23'h00_0000;
      p16_uge_4144 <= 1'h0;
      p16_b_fractionivisor__1 <= 24'h00_0000;
      p16_uge_4152 <= 1'h0;
      p16_uge_4223 <= 1'h0;
      p16_uge_4298 <= 1'h0;
      p16_uge_4364 <= 1'h0;
      p16_uge_4430 <= 1'h0;
      p16_uge_4496 <= 1'h0;
      p16_uge_4562 <= 1'h0;
      p16_uge_4628 <= 1'h0;
      p16_uge_4694 <= 1'h0;
      p16_uge_4760 <= 1'h0;
      p16_uge_4826 <= 1'h0;
      p16_uge_4892 <= 1'h0;
      p16_uge_4958 <= 1'h0;
      p16_uge_5024 <= 1'h0;
      p16_concat_5089 <= 23'h00_0000;
      p16_uge_5090 <= 1'h0;
      p16_bit_slice_4011 <= 1'h0;
      p16_bit_slice_4012 <= 1'h0;
      p16_bit_slice_4013 <= 1'h0;
      p16_bit_slice_4014 <= 1'h0;
      p16_bit_slice_4015 <= 1'h0;
      p16_bit_slice_4017 <= 1'h0;
      p16_bit_slice_4018 <= 1'h0;
      p16_flag_zero <= 1'h0;
      p16_result_sign <= 1'h0;
      p16_result_exp <= 8'h00;
      p17_b_fraction <= 23'h00_0000;
      p17_uge_4144 <= 1'h0;
      p17_b_fractionivisor__1 <= 24'h00_0000;
      p17_uge_4152 <= 1'h0;
      p17_uge_4223 <= 1'h0;
      p17_uge_4298 <= 1'h0;
      p17_uge_4364 <= 1'h0;
      p17_uge_4430 <= 1'h0;
      p17_uge_4496 <= 1'h0;
      p17_uge_4562 <= 1'h0;
      p17_uge_4628 <= 1'h0;
      p17_uge_4694 <= 1'h0;
      p17_uge_4760 <= 1'h0;
      p17_uge_4826 <= 1'h0;
      p17_uge_4892 <= 1'h0;
      p17_uge_4958 <= 1'h0;
      p17_uge_5024 <= 1'h0;
      p17_uge_5090 <= 1'h0;
      p17_concat_5155 <= 23'h00_0000;
      p17_uge_5156 <= 1'h0;
      p17_bit_slice_4012 <= 1'h0;
      p17_bit_slice_4013 <= 1'h0;
      p17_bit_slice_4014 <= 1'h0;
      p17_bit_slice_4015 <= 1'h0;
      p17_bit_slice_4017 <= 1'h0;
      p17_bit_slice_4018 <= 1'h0;
      p17_flag_zero <= 1'h0;
      p17_result_sign <= 1'h0;
      p17_result_exp <= 8'h00;
      p18_b_fraction <= 23'h00_0000;
      p18_uge_4144 <= 1'h0;
      p18_b_fractionivisor__1 <= 24'h00_0000;
      p18_uge_4152 <= 1'h0;
      p18_uge_4223 <= 1'h0;
      p18_uge_4298 <= 1'h0;
      p18_uge_4364 <= 1'h0;
      p18_uge_4430 <= 1'h0;
      p18_uge_4496 <= 1'h0;
      p18_uge_4562 <= 1'h0;
      p18_uge_4628 <= 1'h0;
      p18_uge_4694 <= 1'h0;
      p18_uge_4760 <= 1'h0;
      p18_uge_4826 <= 1'h0;
      p18_uge_4892 <= 1'h0;
      p18_uge_4958 <= 1'h0;
      p18_uge_5024 <= 1'h0;
      p18_uge_5090 <= 1'h0;
      p18_uge_5156 <= 1'h0;
      p18_concat_5221 <= 23'h00_0000;
      p18_uge_5222 <= 1'h0;
      p18_bit_slice_4013 <= 1'h0;
      p18_bit_slice_4014 <= 1'h0;
      p18_bit_slice_4015 <= 1'h0;
      p18_bit_slice_4017 <= 1'h0;
      p18_bit_slice_4018 <= 1'h0;
      p18_flag_zero <= 1'h0;
      p18_result_sign <= 1'h0;
      p18_result_exp <= 8'h00;
      p19_b_fraction <= 23'h00_0000;
      p19_uge_4144 <= 1'h0;
      p19_b_fractionivisor__1 <= 24'h00_0000;
      p19_uge_4152 <= 1'h0;
      p19_uge_4223 <= 1'h0;
      p19_uge_4298 <= 1'h0;
      p19_uge_4364 <= 1'h0;
      p19_uge_4430 <= 1'h0;
      p19_uge_4496 <= 1'h0;
      p19_uge_4562 <= 1'h0;
      p19_uge_4628 <= 1'h0;
      p19_uge_4694 <= 1'h0;
      p19_uge_4760 <= 1'h0;
      p19_uge_4826 <= 1'h0;
      p19_uge_4892 <= 1'h0;
      p19_uge_4958 <= 1'h0;
      p19_uge_5024 <= 1'h0;
      p19_uge_5090 <= 1'h0;
      p19_uge_5156 <= 1'h0;
      p19_uge_5222 <= 1'h0;
      p19_concat_5287 <= 23'h00_0000;
      p19_uge_5288 <= 1'h0;
      p19_bit_slice_4014 <= 1'h0;
      p19_bit_slice_4015 <= 1'h0;
      p19_bit_slice_4017 <= 1'h0;
      p19_bit_slice_4018 <= 1'h0;
      p19_flag_zero <= 1'h0;
      p19_result_sign <= 1'h0;
      p19_result_exp <= 8'h00;
      p20_b_fraction <= 23'h00_0000;
      p20_uge_4144 <= 1'h0;
      p20_b_fractionivisor__1 <= 24'h00_0000;
      p20_uge_4152 <= 1'h0;
      p20_uge_4223 <= 1'h0;
      p20_uge_4298 <= 1'h0;
      p20_uge_4364 <= 1'h0;
      p20_uge_4430 <= 1'h0;
      p20_uge_4496 <= 1'h0;
      p20_uge_4562 <= 1'h0;
      p20_uge_4628 <= 1'h0;
      p20_uge_4694 <= 1'h0;
      p20_uge_4760 <= 1'h0;
      p20_uge_4826 <= 1'h0;
      p20_uge_4892 <= 1'h0;
      p20_uge_4958 <= 1'h0;
      p20_uge_5024 <= 1'h0;
      p20_uge_5090 <= 1'h0;
      p20_uge_5156 <= 1'h0;
      p20_uge_5222 <= 1'h0;
      p20_uge_5288 <= 1'h0;
      p20_concat_5353 <= 23'h00_0000;
      p20_uge_5354 <= 1'h0;
      p20_bit_slice_4015 <= 1'h0;
      p20_bit_slice_4017 <= 1'h0;
      p20_bit_slice_4018 <= 1'h0;
      p20_flag_zero <= 1'h0;
      p20_result_sign <= 1'h0;
      p20_result_exp <= 8'h00;
      p21_b_fraction <= 23'h00_0000;
      p21_uge_4144 <= 1'h0;
      p21_b_fractionivisor__1 <= 24'h00_0000;
      p21_uge_4152 <= 1'h0;
      p21_uge_4223 <= 1'h0;
      p21_uge_4298 <= 1'h0;
      p21_uge_4364 <= 1'h0;
      p21_uge_4430 <= 1'h0;
      p21_uge_4496 <= 1'h0;
      p21_uge_4562 <= 1'h0;
      p21_uge_4628 <= 1'h0;
      p21_uge_4694 <= 1'h0;
      p21_uge_4760 <= 1'h0;
      p21_uge_4826 <= 1'h0;
      p21_uge_4892 <= 1'h0;
      p21_uge_4958 <= 1'h0;
      p21_uge_5024 <= 1'h0;
      p21_uge_5090 <= 1'h0;
      p21_uge_5156 <= 1'h0;
      p21_uge_5222 <= 1'h0;
      p21_uge_5288 <= 1'h0;
      p21_uge_5354 <= 1'h0;
      p21_concat_5419 <= 23'h00_0000;
      p21_uge_5420 <= 1'h0;
      p21_bit_slice_4017 <= 1'h0;
      p21_bit_slice_4018 <= 1'h0;
      p21_flag_zero <= 1'h0;
      p21_result_sign <= 1'h0;
      p21_result_exp <= 8'h00;
      p22_b_fraction <= 23'h00_0000;
      p22_uge_4144 <= 1'h0;
      p22_b_fractionivisor__1 <= 24'h00_0000;
      p22_uge_4152 <= 1'h0;
      p22_uge_4223 <= 1'h0;
      p22_uge_4298 <= 1'h0;
      p22_uge_4364 <= 1'h0;
      p22_uge_4430 <= 1'h0;
      p22_uge_4496 <= 1'h0;
      p22_uge_4562 <= 1'h0;
      p22_uge_4628 <= 1'h0;
      p22_uge_4694 <= 1'h0;
      p22_uge_4760 <= 1'h0;
      p22_uge_4826 <= 1'h0;
      p22_uge_4892 <= 1'h0;
      p22_uge_4958 <= 1'h0;
      p22_uge_5024 <= 1'h0;
      p22_uge_5090 <= 1'h0;
      p22_uge_5156 <= 1'h0;
      p22_uge_5222 <= 1'h0;
      p22_uge_5288 <= 1'h0;
      p22_uge_5354 <= 1'h0;
      p22_uge_5420 <= 1'h0;
      p22_concat_5485 <= 23'h00_0000;
      p22_uge_5486 <= 1'h0;
      p22_bit_slice_4018 <= 1'h0;
      p22_flag_zero <= 1'h0;
      p22_result_sign <= 1'h0;
      p22_result_exp <= 8'h00;
      p23_uge_4144 <= 1'h0;
      p23_uge_4152 <= 1'h0;
      p23_uge_4223 <= 1'h0;
      p23_uge_4298 <= 1'h0;
      p23_uge_4364 <= 1'h0;
      p23_uge_4430 <= 1'h0;
      p23_uge_4496 <= 1'h0;
      p23_uge_4562 <= 1'h0;
      p23_uge_4628 <= 1'h0;
      p23_uge_4694 <= 1'h0;
      p23_uge_4760 <= 1'h0;
      p23_uge_4826 <= 1'h0;
      p23_uge_4892 <= 1'h0;
      p23_uge_4958 <= 1'h0;
      p23_uge_5024 <= 1'h0;
      p23_uge_5090 <= 1'h0;
      p23_uge_5156 <= 1'h0;
      p23_uge_5222 <= 1'h0;
      p23_uge_5288 <= 1'h0;
      p23_uge_5354 <= 1'h0;
      p23_uge_5420 <= 1'h0;
      p23_uge_5486 <= 1'h0;
      p23_flag_zero <= 1'h0;
      p23_q__23_squeezed_portion_0_width_1 <= 1'h0;
      p23_result_sign <= 1'h0;
      p23_result_exp <= 8'h00;
      p0_valid <= 1'h0;
      p1_valid <= 1'h0;
      p2_valid <= 1'h0;
      p3_valid <= 1'h0;
      p4_valid <= 1'h0;
      p5_valid <= 1'h0;
      p6_valid <= 1'h0;
      p7_valid <= 1'h0;
      p8_valid <= 1'h0;
      p9_valid <= 1'h0;
      p10_valid <= 1'h0;
      p11_valid <= 1'h0;
      p12_valid <= 1'h0;
      p13_valid <= 1'h0;
      p14_valid <= 1'h0;
      p15_valid <= 1'h0;
      p16_valid <= 1'h0;
      p17_valid <= 1'h0;
      p18_valid <= 1'h0;
      p19_valid <= 1'h0;
      p20_valid <= 1'h0;
      p21_valid <= 1'h0;
      p22_valid <= 1'h0;
      p23_valid <= 1'h0;
      p24_valid <= 1'h0;
      p25_valid <= 1'h0;
      p26_valid <= 1'h0;
      p27_valid <= 1'h0;
      p28_valid <= 1'h0;
      __xls_float_ips__result_reg <= __xls_float_ips__result_reg_init;
      __xls_float_ips__result_valid_reg <= 1'h0;
    end else begin
      p0_bit_slice_3995 <= p0_data_enable ? bit_slice_3995 : p0_bit_slice_3995;
      p0_bit_slice_3996 <= p0_data_enable ? bit_slice_3996 : p0_bit_slice_3996;
      p0_bit_slice_3997 <= p0_data_enable ? bit_slice_3997 : p0_bit_slice_3997;
      p0_bit_slice_3998 <= p0_data_enable ? bit_slice_3998 : p0_bit_slice_3998;
      p0_bit_slice_3999 <= p0_data_enable ? bit_slice_3999 : p0_bit_slice_3999;
      p0_bit_slice_4000 <= p0_data_enable ? bit_slice_4000 : p0_bit_slice_4000;
      p0_bit_slice_4001 <= p0_data_enable ? bit_slice_4001 : p0_bit_slice_4001;
      p0_bit_slice_4002 <= p0_data_enable ? bit_slice_4002 : p0_bit_slice_4002;
      p0_bit_slice_4003 <= p0_data_enable ? bit_slice_4003 : p0_bit_slice_4003;
      p0_bit_slice_4004 <= p0_data_enable ? bit_slice_4004 : p0_bit_slice_4004;
      p0_bit_slice_4005 <= p0_data_enable ? bit_slice_4005 : p0_bit_slice_4005;
      p0_bit_slice_4006 <= p0_data_enable ? bit_slice_4006 : p0_bit_slice_4006;
      p0_bit_slice_4007 <= p0_data_enable ? bit_slice_4007 : p0_bit_slice_4007;
      p0_bit_slice_4008 <= p0_data_enable ? bit_slice_4008 : p0_bit_slice_4008;
      p0_bit_slice_4009 <= p0_data_enable ? bit_slice_4009 : p0_bit_slice_4009;
      p0_bit_slice_4010 <= p0_data_enable ? bit_slice_4010 : p0_bit_slice_4010;
      p0_bit_slice_4011 <= p0_data_enable ? bit_slice_4011 : p0_bit_slice_4011;
      p0_bit_slice_4012 <= p0_data_enable ? bit_slice_4012 : p0_bit_slice_4012;
      p0_bit_slice_4013 <= p0_data_enable ? bit_slice_4013 : p0_bit_slice_4013;
      p0_bit_slice_4014 <= p0_data_enable ? bit_slice_4014 : p0_bit_slice_4014;
      p0_bit_slice_4015 <= p0_data_enable ? bit_slice_4015 : p0_bit_slice_4015;
      p0_a_bexp <= p0_data_enable ? a_bexp : p0_a_bexp;
      p0_bit_slice_4017 <= p0_data_enable ? bit_slice_4017 : p0_bit_slice_4017;
      p0_bit_slice_4018 <= p0_data_enable ? bit_slice_4018 : p0_bit_slice_4018;
      p0_a_sign <= p0_data_enable ? a_sign : p0_a_sign;
      p1_concat_4081 <= p1_data_enable ? concat_4081 : p1_concat_4081;
      p1_b_fraction <= p1_data_enable ? b_fraction : p1_b_fraction;
      p1_bit_slice_3996 <= p1_data_enable ? p0_bit_slice_3996 : p1_bit_slice_3996;
      p1_bit_slice_3997 <= p1_data_enable ? p0_bit_slice_3997 : p1_bit_slice_3997;
      p1_bit_slice_3998 <= p1_data_enable ? p0_bit_slice_3998 : p1_bit_slice_3998;
      p1_bit_slice_3999 <= p1_data_enable ? p0_bit_slice_3999 : p1_bit_slice_3999;
      p1_bit_slice_4000 <= p1_data_enable ? p0_bit_slice_4000 : p1_bit_slice_4000;
      p1_bit_slice_4001 <= p1_data_enable ? p0_bit_slice_4001 : p1_bit_slice_4001;
      p1_bit_slice_4002 <= p1_data_enable ? p0_bit_slice_4002 : p1_bit_slice_4002;
      p1_bit_slice_4003 <= p1_data_enable ? p0_bit_slice_4003 : p1_bit_slice_4003;
      p1_bit_slice_4004 <= p1_data_enable ? p0_bit_slice_4004 : p1_bit_slice_4004;
      p1_bit_slice_4005 <= p1_data_enable ? p0_bit_slice_4005 : p1_bit_slice_4005;
      p1_bit_slice_4006 <= p1_data_enable ? p0_bit_slice_4006 : p1_bit_slice_4006;
      p1_bit_slice_4007 <= p1_data_enable ? p0_bit_slice_4007 : p1_bit_slice_4007;
      p1_bit_slice_4008 <= p1_data_enable ? p0_bit_slice_4008 : p1_bit_slice_4008;
      p1_bit_slice_4009 <= p1_data_enable ? p0_bit_slice_4009 : p1_bit_slice_4009;
      p1_bit_slice_4010 <= p1_data_enable ? p0_bit_slice_4010 : p1_bit_slice_4010;
      p1_bit_slice_4011 <= p1_data_enable ? p0_bit_slice_4011 : p1_bit_slice_4011;
      p1_bit_slice_4012 <= p1_data_enable ? p0_bit_slice_4012 : p1_bit_slice_4012;
      p1_bit_slice_4013 <= p1_data_enable ? p0_bit_slice_4013 : p1_bit_slice_4013;
      p1_bit_slice_4014 <= p1_data_enable ? p0_bit_slice_4014 : p1_bit_slice_4014;
      p1_bit_slice_4015 <= p1_data_enable ? p0_bit_slice_4015 : p1_bit_slice_4015;
      p1_a_bexp <= p1_data_enable ? p0_a_bexp : p1_a_bexp;
      p1_b_bexp <= p1_data_enable ? b_bexp : p1_b_bexp;
      p1_bit_slice_4017 <= p1_data_enable ? p0_bit_slice_4017 : p1_bit_slice_4017;
      p1_bit_slice_4018 <= p1_data_enable ? p0_bit_slice_4018 : p1_bit_slice_4018;
      p1_result_sign <= p1_data_enable ? result_sign : p1_result_sign;
      p2_b_fraction <= p2_data_enable ? p1_b_fraction : p2_b_fraction;
      p2_uge_4144 <= p2_data_enable ? uge_4144 : p2_uge_4144;
      p2_b_fractionivisor__1 <= p2_data_enable ? b_fractionivisor__1 : p2_b_fractionivisor__1;
      p2_concat_4151 <= p2_data_enable ? concat_4151 : p2_concat_4151;
      p2_uge_4152 <= p2_data_enable ? uge_4152 : p2_uge_4152;
      p2_bit_slice_3997 <= p2_data_enable ? p1_bit_slice_3997 : p2_bit_slice_3997;
      p2_bit_slice_3998 <= p2_data_enable ? p1_bit_slice_3998 : p2_bit_slice_3998;
      p2_bit_slice_3999 <= p2_data_enable ? p1_bit_slice_3999 : p2_bit_slice_3999;
      p2_bit_slice_4000 <= p2_data_enable ? p1_bit_slice_4000 : p2_bit_slice_4000;
      p2_bit_slice_4001 <= p2_data_enable ? p1_bit_slice_4001 : p2_bit_slice_4001;
      p2_bit_slice_4002 <= p2_data_enable ? p1_bit_slice_4002 : p2_bit_slice_4002;
      p2_bit_slice_4003 <= p2_data_enable ? p1_bit_slice_4003 : p2_bit_slice_4003;
      p2_bit_slice_4004 <= p2_data_enable ? p1_bit_slice_4004 : p2_bit_slice_4004;
      p2_bit_slice_4005 <= p2_data_enable ? p1_bit_slice_4005 : p2_bit_slice_4005;
      p2_bit_slice_4006 <= p2_data_enable ? p1_bit_slice_4006 : p2_bit_slice_4006;
      p2_bit_slice_4007 <= p2_data_enable ? p1_bit_slice_4007 : p2_bit_slice_4007;
      p2_bit_slice_4008 <= p2_data_enable ? p1_bit_slice_4008 : p2_bit_slice_4008;
      p2_bit_slice_4009 <= p2_data_enable ? p1_bit_slice_4009 : p2_bit_slice_4009;
      p2_bit_slice_4010 <= p2_data_enable ? p1_bit_slice_4010 : p2_bit_slice_4010;
      p2_bit_slice_4011 <= p2_data_enable ? p1_bit_slice_4011 : p2_bit_slice_4011;
      p2_bit_slice_4012 <= p2_data_enable ? p1_bit_slice_4012 : p2_bit_slice_4012;
      p2_bit_slice_4013 <= p2_data_enable ? p1_bit_slice_4013 : p2_bit_slice_4013;
      p2_bit_slice_4014 <= p2_data_enable ? p1_bit_slice_4014 : p2_bit_slice_4014;
      p2_bit_slice_4015 <= p2_data_enable ? p1_bit_slice_4015 : p2_bit_slice_4015;
      p2_bit_slice_4017 <= p2_data_enable ? p1_bit_slice_4017 : p2_bit_slice_4017;
      p2_signed_exp_s9 <= p2_data_enable ? signed_exp_s9 : p2_signed_exp_s9;
      p2_bit_slice_4018 <= p2_data_enable ? p1_bit_slice_4018 : p2_bit_slice_4018;
      p2_result_sign <= p2_data_enable ? p1_result_sign : p2_result_sign;
      p3_b_fraction <= p3_data_enable ? p2_b_fraction : p3_b_fraction;
      p3_uge_4144 <= p3_data_enable ? p2_uge_4144 : p3_uge_4144;
      p3_b_fractionivisor__1 <= p3_data_enable ? p2_b_fractionivisor__1 : p3_b_fractionivisor__1;
      p3_uge_4152 <= p3_data_enable ? p2_uge_4152 : p3_uge_4152;
      p3_concat_4222 <= p3_data_enable ? concat_4222 : p3_concat_4222;
      p3_uge_4223 <= p3_data_enable ? uge_4223 : p3_uge_4223;
      p3_bit_slice_3998 <= p3_data_enable ? p2_bit_slice_3998 : p3_bit_slice_3998;
      p3_bit_slice_3999 <= p3_data_enable ? p2_bit_slice_3999 : p3_bit_slice_3999;
      p3_bit_slice_4000 <= p3_data_enable ? p2_bit_slice_4000 : p3_bit_slice_4000;
      p3_bit_slice_4001 <= p3_data_enable ? p2_bit_slice_4001 : p3_bit_slice_4001;
      p3_bit_slice_4002 <= p3_data_enable ? p2_bit_slice_4002 : p3_bit_slice_4002;
      p3_bit_slice_4003 <= p3_data_enable ? p2_bit_slice_4003 : p3_bit_slice_4003;
      p3_bit_slice_4004 <= p3_data_enable ? p2_bit_slice_4004 : p3_bit_slice_4004;
      p3_bit_slice_4005 <= p3_data_enable ? p2_bit_slice_4005 : p3_bit_slice_4005;
      p3_bit_slice_4006 <= p3_data_enable ? p2_bit_slice_4006 : p3_bit_slice_4006;
      p3_bit_slice_4007 <= p3_data_enable ? p2_bit_slice_4007 : p3_bit_slice_4007;
      p3_bit_slice_4008 <= p3_data_enable ? p2_bit_slice_4008 : p3_bit_slice_4008;
      p3_bit_slice_4009 <= p3_data_enable ? p2_bit_slice_4009 : p3_bit_slice_4009;
      p3_bit_slice_4010 <= p3_data_enable ? p2_bit_slice_4010 : p3_bit_slice_4010;
      p3_bit_slice_4011 <= p3_data_enable ? p2_bit_slice_4011 : p3_bit_slice_4011;
      p3_bit_slice_4012 <= p3_data_enable ? p2_bit_slice_4012 : p3_bit_slice_4012;
      p3_bit_slice_4013 <= p3_data_enable ? p2_bit_slice_4013 : p3_bit_slice_4013;
      p3_bit_slice_4014 <= p3_data_enable ? p2_bit_slice_4014 : p3_bit_slice_4014;
      p3_bit_slice_4015 <= p3_data_enable ? p2_bit_slice_4015 : p3_bit_slice_4015;
      p3_bit_slice_4017 <= p3_data_enable ? p2_bit_slice_4017 : p3_bit_slice_4017;
      p3_bit_slice_4018 <= p3_data_enable ? p2_bit_slice_4018 : p3_bit_slice_4018;
      p3_flag_zero <= p3_data_enable ? flag_zero : p3_flag_zero;
      p3_result_sign <= p3_data_enable ? p2_result_sign : p3_result_sign;
      p3_result_exp <= p3_data_enable ? result_exp : p3_result_exp;
      p4_b_fraction <= p4_data_enable ? p3_b_fraction : p4_b_fraction;
      p4_uge_4144 <= p4_data_enable ? p3_uge_4144 : p4_uge_4144;
      p4_b_fractionivisor__1 <= p4_data_enable ? p3_b_fractionivisor__1 : p4_b_fractionivisor__1;
      p4_uge_4152 <= p4_data_enable ? p3_uge_4152 : p4_uge_4152;
      p4_uge_4223 <= p4_data_enable ? p3_uge_4223 : p4_uge_4223;
      p4_concat_4297 <= p4_data_enable ? concat_4297 : p4_concat_4297;
      p4_uge_4298 <= p4_data_enable ? uge_4298 : p4_uge_4298;
      p4_bit_slice_3999 <= p4_data_enable ? p3_bit_slice_3999 : p4_bit_slice_3999;
      p4_bit_slice_4000 <= p4_data_enable ? p3_bit_slice_4000 : p4_bit_slice_4000;
      p4_bit_slice_4001 <= p4_data_enable ? p3_bit_slice_4001 : p4_bit_slice_4001;
      p4_bit_slice_4002 <= p4_data_enable ? p3_bit_slice_4002 : p4_bit_slice_4002;
      p4_bit_slice_4003 <= p4_data_enable ? p3_bit_slice_4003 : p4_bit_slice_4003;
      p4_bit_slice_4004 <= p4_data_enable ? p3_bit_slice_4004 : p4_bit_slice_4004;
      p4_bit_slice_4005 <= p4_data_enable ? p3_bit_slice_4005 : p4_bit_slice_4005;
      p4_bit_slice_4006 <= p4_data_enable ? p3_bit_slice_4006 : p4_bit_slice_4006;
      p4_bit_slice_4007 <= p4_data_enable ? p3_bit_slice_4007 : p4_bit_slice_4007;
      p4_bit_slice_4008 <= p4_data_enable ? p3_bit_slice_4008 : p4_bit_slice_4008;
      p4_bit_slice_4009 <= p4_data_enable ? p3_bit_slice_4009 : p4_bit_slice_4009;
      p4_bit_slice_4010 <= p4_data_enable ? p3_bit_slice_4010 : p4_bit_slice_4010;
      p4_bit_slice_4011 <= p4_data_enable ? p3_bit_slice_4011 : p4_bit_slice_4011;
      p4_bit_slice_4012 <= p4_data_enable ? p3_bit_slice_4012 : p4_bit_slice_4012;
      p4_bit_slice_4013 <= p4_data_enable ? p3_bit_slice_4013 : p4_bit_slice_4013;
      p4_bit_slice_4014 <= p4_data_enable ? p3_bit_slice_4014 : p4_bit_slice_4014;
      p4_bit_slice_4015 <= p4_data_enable ? p3_bit_slice_4015 : p4_bit_slice_4015;
      p4_bit_slice_4017 <= p4_data_enable ? p3_bit_slice_4017 : p4_bit_slice_4017;
      p4_bit_slice_4018 <= p4_data_enable ? p3_bit_slice_4018 : p4_bit_slice_4018;
      p4_flag_zero <= p4_data_enable ? p3_flag_zero : p4_flag_zero;
      p4_result_sign <= p4_data_enable ? p3_result_sign : p4_result_sign;
      p4_result_exp <= p4_data_enable ? p3_result_exp : p4_result_exp;
      p5_b_fraction <= p5_data_enable ? p4_b_fraction : p5_b_fraction;
      p5_uge_4144 <= p5_data_enable ? p4_uge_4144 : p5_uge_4144;
      p5_b_fractionivisor__1 <= p5_data_enable ? p4_b_fractionivisor__1 : p5_b_fractionivisor__1;
      p5_uge_4152 <= p5_data_enable ? p4_uge_4152 : p5_uge_4152;
      p5_uge_4223 <= p5_data_enable ? p4_uge_4223 : p5_uge_4223;
      p5_uge_4298 <= p5_data_enable ? p4_uge_4298 : p5_uge_4298;
      p5_concat_4363 <= p5_data_enable ? concat_4363 : p5_concat_4363;
      p5_uge_4364 <= p5_data_enable ? uge_4364 : p5_uge_4364;
      p5_bit_slice_4000 <= p5_data_enable ? p4_bit_slice_4000 : p5_bit_slice_4000;
      p5_bit_slice_4001 <= p5_data_enable ? p4_bit_slice_4001 : p5_bit_slice_4001;
      p5_bit_slice_4002 <= p5_data_enable ? p4_bit_slice_4002 : p5_bit_slice_4002;
      p5_bit_slice_4003 <= p5_data_enable ? p4_bit_slice_4003 : p5_bit_slice_4003;
      p5_bit_slice_4004 <= p5_data_enable ? p4_bit_slice_4004 : p5_bit_slice_4004;
      p5_bit_slice_4005 <= p5_data_enable ? p4_bit_slice_4005 : p5_bit_slice_4005;
      p5_bit_slice_4006 <= p5_data_enable ? p4_bit_slice_4006 : p5_bit_slice_4006;
      p5_bit_slice_4007 <= p5_data_enable ? p4_bit_slice_4007 : p5_bit_slice_4007;
      p5_bit_slice_4008 <= p5_data_enable ? p4_bit_slice_4008 : p5_bit_slice_4008;
      p5_bit_slice_4009 <= p5_data_enable ? p4_bit_slice_4009 : p5_bit_slice_4009;
      p5_bit_slice_4010 <= p5_data_enable ? p4_bit_slice_4010 : p5_bit_slice_4010;
      p5_bit_slice_4011 <= p5_data_enable ? p4_bit_slice_4011 : p5_bit_slice_4011;
      p5_bit_slice_4012 <= p5_data_enable ? p4_bit_slice_4012 : p5_bit_slice_4012;
      p5_bit_slice_4013 <= p5_data_enable ? p4_bit_slice_4013 : p5_bit_slice_4013;
      p5_bit_slice_4014 <= p5_data_enable ? p4_bit_slice_4014 : p5_bit_slice_4014;
      p5_bit_slice_4015 <= p5_data_enable ? p4_bit_slice_4015 : p5_bit_slice_4015;
      p5_bit_slice_4017 <= p5_data_enable ? p4_bit_slice_4017 : p5_bit_slice_4017;
      p5_bit_slice_4018 <= p5_data_enable ? p4_bit_slice_4018 : p5_bit_slice_4018;
      p5_flag_zero <= p5_data_enable ? p4_flag_zero : p5_flag_zero;
      p5_result_sign <= p5_data_enable ? p4_result_sign : p5_result_sign;
      p5_result_exp <= p5_data_enable ? p4_result_exp : p5_result_exp;
      p6_b_fraction <= p6_data_enable ? p5_b_fraction : p6_b_fraction;
      p6_uge_4144 <= p6_data_enable ? p5_uge_4144 : p6_uge_4144;
      p6_b_fractionivisor__1 <= p6_data_enable ? p5_b_fractionivisor__1 : p6_b_fractionivisor__1;
      p6_uge_4152 <= p6_data_enable ? p5_uge_4152 : p6_uge_4152;
      p6_uge_4223 <= p6_data_enable ? p5_uge_4223 : p6_uge_4223;
      p6_uge_4298 <= p6_data_enable ? p5_uge_4298 : p6_uge_4298;
      p6_uge_4364 <= p6_data_enable ? p5_uge_4364 : p6_uge_4364;
      p6_concat_4429 <= p6_data_enable ? concat_4429 : p6_concat_4429;
      p6_uge_4430 <= p6_data_enable ? uge_4430 : p6_uge_4430;
      p6_bit_slice_4001 <= p6_data_enable ? p5_bit_slice_4001 : p6_bit_slice_4001;
      p6_bit_slice_4002 <= p6_data_enable ? p5_bit_slice_4002 : p6_bit_slice_4002;
      p6_bit_slice_4003 <= p6_data_enable ? p5_bit_slice_4003 : p6_bit_slice_4003;
      p6_bit_slice_4004 <= p6_data_enable ? p5_bit_slice_4004 : p6_bit_slice_4004;
      p6_bit_slice_4005 <= p6_data_enable ? p5_bit_slice_4005 : p6_bit_slice_4005;
      p6_bit_slice_4006 <= p6_data_enable ? p5_bit_slice_4006 : p6_bit_slice_4006;
      p6_bit_slice_4007 <= p6_data_enable ? p5_bit_slice_4007 : p6_bit_slice_4007;
      p6_bit_slice_4008 <= p6_data_enable ? p5_bit_slice_4008 : p6_bit_slice_4008;
      p6_bit_slice_4009 <= p6_data_enable ? p5_bit_slice_4009 : p6_bit_slice_4009;
      p6_bit_slice_4010 <= p6_data_enable ? p5_bit_slice_4010 : p6_bit_slice_4010;
      p6_bit_slice_4011 <= p6_data_enable ? p5_bit_slice_4011 : p6_bit_slice_4011;
      p6_bit_slice_4012 <= p6_data_enable ? p5_bit_slice_4012 : p6_bit_slice_4012;
      p6_bit_slice_4013 <= p6_data_enable ? p5_bit_slice_4013 : p6_bit_slice_4013;
      p6_bit_slice_4014 <= p6_data_enable ? p5_bit_slice_4014 : p6_bit_slice_4014;
      p6_bit_slice_4015 <= p6_data_enable ? p5_bit_slice_4015 : p6_bit_slice_4015;
      p6_bit_slice_4017 <= p6_data_enable ? p5_bit_slice_4017 : p6_bit_slice_4017;
      p6_bit_slice_4018 <= p6_data_enable ? p5_bit_slice_4018 : p6_bit_slice_4018;
      p6_flag_zero <= p6_data_enable ? p5_flag_zero : p6_flag_zero;
      p6_result_sign <= p6_data_enable ? p5_result_sign : p6_result_sign;
      p6_result_exp <= p6_data_enable ? p5_result_exp : p6_result_exp;
      p7_b_fraction <= p7_data_enable ? p6_b_fraction : p7_b_fraction;
      p7_uge_4144 <= p7_data_enable ? p6_uge_4144 : p7_uge_4144;
      p7_b_fractionivisor__1 <= p7_data_enable ? p6_b_fractionivisor__1 : p7_b_fractionivisor__1;
      p7_uge_4152 <= p7_data_enable ? p6_uge_4152 : p7_uge_4152;
      p7_uge_4223 <= p7_data_enable ? p6_uge_4223 : p7_uge_4223;
      p7_uge_4298 <= p7_data_enable ? p6_uge_4298 : p7_uge_4298;
      p7_uge_4364 <= p7_data_enable ? p6_uge_4364 : p7_uge_4364;
      p7_uge_4430 <= p7_data_enable ? p6_uge_4430 : p7_uge_4430;
      p7_concat_4495 <= p7_data_enable ? concat_4495 : p7_concat_4495;
      p7_uge_4496 <= p7_data_enable ? uge_4496 : p7_uge_4496;
      p7_bit_slice_4002 <= p7_data_enable ? p6_bit_slice_4002 : p7_bit_slice_4002;
      p7_bit_slice_4003 <= p7_data_enable ? p6_bit_slice_4003 : p7_bit_slice_4003;
      p7_bit_slice_4004 <= p7_data_enable ? p6_bit_slice_4004 : p7_bit_slice_4004;
      p7_bit_slice_4005 <= p7_data_enable ? p6_bit_slice_4005 : p7_bit_slice_4005;
      p7_bit_slice_4006 <= p7_data_enable ? p6_bit_slice_4006 : p7_bit_slice_4006;
      p7_bit_slice_4007 <= p7_data_enable ? p6_bit_slice_4007 : p7_bit_slice_4007;
      p7_bit_slice_4008 <= p7_data_enable ? p6_bit_slice_4008 : p7_bit_slice_4008;
      p7_bit_slice_4009 <= p7_data_enable ? p6_bit_slice_4009 : p7_bit_slice_4009;
      p7_bit_slice_4010 <= p7_data_enable ? p6_bit_slice_4010 : p7_bit_slice_4010;
      p7_bit_slice_4011 <= p7_data_enable ? p6_bit_slice_4011 : p7_bit_slice_4011;
      p7_bit_slice_4012 <= p7_data_enable ? p6_bit_slice_4012 : p7_bit_slice_4012;
      p7_bit_slice_4013 <= p7_data_enable ? p6_bit_slice_4013 : p7_bit_slice_4013;
      p7_bit_slice_4014 <= p7_data_enable ? p6_bit_slice_4014 : p7_bit_slice_4014;
      p7_bit_slice_4015 <= p7_data_enable ? p6_bit_slice_4015 : p7_bit_slice_4015;
      p7_bit_slice_4017 <= p7_data_enable ? p6_bit_slice_4017 : p7_bit_slice_4017;
      p7_bit_slice_4018 <= p7_data_enable ? p6_bit_slice_4018 : p7_bit_slice_4018;
      p7_flag_zero <= p7_data_enable ? p6_flag_zero : p7_flag_zero;
      p7_result_sign <= p7_data_enable ? p6_result_sign : p7_result_sign;
      p7_result_exp <= p7_data_enable ? p6_result_exp : p7_result_exp;
      p8_b_fraction <= p8_data_enable ? p7_b_fraction : p8_b_fraction;
      p8_uge_4144 <= p8_data_enable ? p7_uge_4144 : p8_uge_4144;
      p8_b_fractionivisor__1 <= p8_data_enable ? p7_b_fractionivisor__1 : p8_b_fractionivisor__1;
      p8_uge_4152 <= p8_data_enable ? p7_uge_4152 : p8_uge_4152;
      p8_uge_4223 <= p8_data_enable ? p7_uge_4223 : p8_uge_4223;
      p8_uge_4298 <= p8_data_enable ? p7_uge_4298 : p8_uge_4298;
      p8_uge_4364 <= p8_data_enable ? p7_uge_4364 : p8_uge_4364;
      p8_uge_4430 <= p8_data_enable ? p7_uge_4430 : p8_uge_4430;
      p8_uge_4496 <= p8_data_enable ? p7_uge_4496 : p8_uge_4496;
      p8_concat_4561 <= p8_data_enable ? concat_4561 : p8_concat_4561;
      p8_uge_4562 <= p8_data_enable ? uge_4562 : p8_uge_4562;
      p8_bit_slice_4003 <= p8_data_enable ? p7_bit_slice_4003 : p8_bit_slice_4003;
      p8_bit_slice_4004 <= p8_data_enable ? p7_bit_slice_4004 : p8_bit_slice_4004;
      p8_bit_slice_4005 <= p8_data_enable ? p7_bit_slice_4005 : p8_bit_slice_4005;
      p8_bit_slice_4006 <= p8_data_enable ? p7_bit_slice_4006 : p8_bit_slice_4006;
      p8_bit_slice_4007 <= p8_data_enable ? p7_bit_slice_4007 : p8_bit_slice_4007;
      p8_bit_slice_4008 <= p8_data_enable ? p7_bit_slice_4008 : p8_bit_slice_4008;
      p8_bit_slice_4009 <= p8_data_enable ? p7_bit_slice_4009 : p8_bit_slice_4009;
      p8_bit_slice_4010 <= p8_data_enable ? p7_bit_slice_4010 : p8_bit_slice_4010;
      p8_bit_slice_4011 <= p8_data_enable ? p7_bit_slice_4011 : p8_bit_slice_4011;
      p8_bit_slice_4012 <= p8_data_enable ? p7_bit_slice_4012 : p8_bit_slice_4012;
      p8_bit_slice_4013 <= p8_data_enable ? p7_bit_slice_4013 : p8_bit_slice_4013;
      p8_bit_slice_4014 <= p8_data_enable ? p7_bit_slice_4014 : p8_bit_slice_4014;
      p8_bit_slice_4015 <= p8_data_enable ? p7_bit_slice_4015 : p8_bit_slice_4015;
      p8_bit_slice_4017 <= p8_data_enable ? p7_bit_slice_4017 : p8_bit_slice_4017;
      p8_bit_slice_4018 <= p8_data_enable ? p7_bit_slice_4018 : p8_bit_slice_4018;
      p8_flag_zero <= p8_data_enable ? p7_flag_zero : p8_flag_zero;
      p8_result_sign <= p8_data_enable ? p7_result_sign : p8_result_sign;
      p8_result_exp <= p8_data_enable ? p7_result_exp : p8_result_exp;
      p9_b_fraction <= p9_data_enable ? p8_b_fraction : p9_b_fraction;
      p9_uge_4144 <= p9_data_enable ? p8_uge_4144 : p9_uge_4144;
      p9_b_fractionivisor__1 <= p9_data_enable ? p8_b_fractionivisor__1 : p9_b_fractionivisor__1;
      p9_uge_4152 <= p9_data_enable ? p8_uge_4152 : p9_uge_4152;
      p9_uge_4223 <= p9_data_enable ? p8_uge_4223 : p9_uge_4223;
      p9_uge_4298 <= p9_data_enable ? p8_uge_4298 : p9_uge_4298;
      p9_uge_4364 <= p9_data_enable ? p8_uge_4364 : p9_uge_4364;
      p9_uge_4430 <= p9_data_enable ? p8_uge_4430 : p9_uge_4430;
      p9_uge_4496 <= p9_data_enable ? p8_uge_4496 : p9_uge_4496;
      p9_uge_4562 <= p9_data_enable ? p8_uge_4562 : p9_uge_4562;
      p9_concat_4627 <= p9_data_enable ? concat_4627 : p9_concat_4627;
      p9_uge_4628 <= p9_data_enable ? uge_4628 : p9_uge_4628;
      p9_bit_slice_4004 <= p9_data_enable ? p8_bit_slice_4004 : p9_bit_slice_4004;
      p9_bit_slice_4005 <= p9_data_enable ? p8_bit_slice_4005 : p9_bit_slice_4005;
      p9_bit_slice_4006 <= p9_data_enable ? p8_bit_slice_4006 : p9_bit_slice_4006;
      p9_bit_slice_4007 <= p9_data_enable ? p8_bit_slice_4007 : p9_bit_slice_4007;
      p9_bit_slice_4008 <= p9_data_enable ? p8_bit_slice_4008 : p9_bit_slice_4008;
      p9_bit_slice_4009 <= p9_data_enable ? p8_bit_slice_4009 : p9_bit_slice_4009;
      p9_bit_slice_4010 <= p9_data_enable ? p8_bit_slice_4010 : p9_bit_slice_4010;
      p9_bit_slice_4011 <= p9_data_enable ? p8_bit_slice_4011 : p9_bit_slice_4011;
      p9_bit_slice_4012 <= p9_data_enable ? p8_bit_slice_4012 : p9_bit_slice_4012;
      p9_bit_slice_4013 <= p9_data_enable ? p8_bit_slice_4013 : p9_bit_slice_4013;
      p9_bit_slice_4014 <= p9_data_enable ? p8_bit_slice_4014 : p9_bit_slice_4014;
      p9_bit_slice_4015 <= p9_data_enable ? p8_bit_slice_4015 : p9_bit_slice_4015;
      p9_bit_slice_4017 <= p9_data_enable ? p8_bit_slice_4017 : p9_bit_slice_4017;
      p9_bit_slice_4018 <= p9_data_enable ? p8_bit_slice_4018 : p9_bit_slice_4018;
      p9_flag_zero <= p9_data_enable ? p8_flag_zero : p9_flag_zero;
      p9_result_sign <= p9_data_enable ? p8_result_sign : p9_result_sign;
      p9_result_exp <= p9_data_enable ? p8_result_exp : p9_result_exp;
      p10_b_fraction <= p10_data_enable ? p9_b_fraction : p10_b_fraction;
      p10_uge_4144 <= p10_data_enable ? p9_uge_4144 : p10_uge_4144;
      p10_b_fractionivisor__1 <= p10_data_enable ? p9_b_fractionivisor__1 : p10_b_fractionivisor__1;
      p10_uge_4152 <= p10_data_enable ? p9_uge_4152 : p10_uge_4152;
      p10_uge_4223 <= p10_data_enable ? p9_uge_4223 : p10_uge_4223;
      p10_uge_4298 <= p10_data_enable ? p9_uge_4298 : p10_uge_4298;
      p10_uge_4364 <= p10_data_enable ? p9_uge_4364 : p10_uge_4364;
      p10_uge_4430 <= p10_data_enable ? p9_uge_4430 : p10_uge_4430;
      p10_uge_4496 <= p10_data_enable ? p9_uge_4496 : p10_uge_4496;
      p10_uge_4562 <= p10_data_enable ? p9_uge_4562 : p10_uge_4562;
      p10_uge_4628 <= p10_data_enable ? p9_uge_4628 : p10_uge_4628;
      p10_concat_4693 <= p10_data_enable ? concat_4693 : p10_concat_4693;
      p10_uge_4694 <= p10_data_enable ? uge_4694 : p10_uge_4694;
      p10_bit_slice_4005 <= p10_data_enable ? p9_bit_slice_4005 : p10_bit_slice_4005;
      p10_bit_slice_4006 <= p10_data_enable ? p9_bit_slice_4006 : p10_bit_slice_4006;
      p10_bit_slice_4007 <= p10_data_enable ? p9_bit_slice_4007 : p10_bit_slice_4007;
      p10_bit_slice_4008 <= p10_data_enable ? p9_bit_slice_4008 : p10_bit_slice_4008;
      p10_bit_slice_4009 <= p10_data_enable ? p9_bit_slice_4009 : p10_bit_slice_4009;
      p10_bit_slice_4010 <= p10_data_enable ? p9_bit_slice_4010 : p10_bit_slice_4010;
      p10_bit_slice_4011 <= p10_data_enable ? p9_bit_slice_4011 : p10_bit_slice_4011;
      p10_bit_slice_4012 <= p10_data_enable ? p9_bit_slice_4012 : p10_bit_slice_4012;
      p10_bit_slice_4013 <= p10_data_enable ? p9_bit_slice_4013 : p10_bit_slice_4013;
      p10_bit_slice_4014 <= p10_data_enable ? p9_bit_slice_4014 : p10_bit_slice_4014;
      p10_bit_slice_4015 <= p10_data_enable ? p9_bit_slice_4015 : p10_bit_slice_4015;
      p10_bit_slice_4017 <= p10_data_enable ? p9_bit_slice_4017 : p10_bit_slice_4017;
      p10_bit_slice_4018 <= p10_data_enable ? p9_bit_slice_4018 : p10_bit_slice_4018;
      p10_flag_zero <= p10_data_enable ? p9_flag_zero : p10_flag_zero;
      p10_result_sign <= p10_data_enable ? p9_result_sign : p10_result_sign;
      p10_result_exp <= p10_data_enable ? p9_result_exp : p10_result_exp;
      p11_b_fraction <= p11_data_enable ? p10_b_fraction : p11_b_fraction;
      p11_uge_4144 <= p11_data_enable ? p10_uge_4144 : p11_uge_4144;
      p11_b_fractionivisor__1 <= p11_data_enable ? p10_b_fractionivisor__1 : p11_b_fractionivisor__1;
      p11_uge_4152 <= p11_data_enable ? p10_uge_4152 : p11_uge_4152;
      p11_uge_4223 <= p11_data_enable ? p10_uge_4223 : p11_uge_4223;
      p11_uge_4298 <= p11_data_enable ? p10_uge_4298 : p11_uge_4298;
      p11_uge_4364 <= p11_data_enable ? p10_uge_4364 : p11_uge_4364;
      p11_uge_4430 <= p11_data_enable ? p10_uge_4430 : p11_uge_4430;
      p11_uge_4496 <= p11_data_enable ? p10_uge_4496 : p11_uge_4496;
      p11_uge_4562 <= p11_data_enable ? p10_uge_4562 : p11_uge_4562;
      p11_uge_4628 <= p11_data_enable ? p10_uge_4628 : p11_uge_4628;
      p11_uge_4694 <= p11_data_enable ? p10_uge_4694 : p11_uge_4694;
      p11_concat_4759 <= p11_data_enable ? concat_4759 : p11_concat_4759;
      p11_uge_4760 <= p11_data_enable ? uge_4760 : p11_uge_4760;
      p11_bit_slice_4006 <= p11_data_enable ? p10_bit_slice_4006 : p11_bit_slice_4006;
      p11_bit_slice_4007 <= p11_data_enable ? p10_bit_slice_4007 : p11_bit_slice_4007;
      p11_bit_slice_4008 <= p11_data_enable ? p10_bit_slice_4008 : p11_bit_slice_4008;
      p11_bit_slice_4009 <= p11_data_enable ? p10_bit_slice_4009 : p11_bit_slice_4009;
      p11_bit_slice_4010 <= p11_data_enable ? p10_bit_slice_4010 : p11_bit_slice_4010;
      p11_bit_slice_4011 <= p11_data_enable ? p10_bit_slice_4011 : p11_bit_slice_4011;
      p11_bit_slice_4012 <= p11_data_enable ? p10_bit_slice_4012 : p11_bit_slice_4012;
      p11_bit_slice_4013 <= p11_data_enable ? p10_bit_slice_4013 : p11_bit_slice_4013;
      p11_bit_slice_4014 <= p11_data_enable ? p10_bit_slice_4014 : p11_bit_slice_4014;
      p11_bit_slice_4015 <= p11_data_enable ? p10_bit_slice_4015 : p11_bit_slice_4015;
      p11_bit_slice_4017 <= p11_data_enable ? p10_bit_slice_4017 : p11_bit_slice_4017;
      p11_bit_slice_4018 <= p11_data_enable ? p10_bit_slice_4018 : p11_bit_slice_4018;
      p11_flag_zero <= p11_data_enable ? p10_flag_zero : p11_flag_zero;
      p11_result_sign <= p11_data_enable ? p10_result_sign : p11_result_sign;
      p11_result_exp <= p11_data_enable ? p10_result_exp : p11_result_exp;
      p12_b_fraction <= p12_data_enable ? p11_b_fraction : p12_b_fraction;
      p12_uge_4144 <= p12_data_enable ? p11_uge_4144 : p12_uge_4144;
      p12_b_fractionivisor__1 <= p12_data_enable ? p11_b_fractionivisor__1 : p12_b_fractionivisor__1;
      p12_uge_4152 <= p12_data_enable ? p11_uge_4152 : p12_uge_4152;
      p12_uge_4223 <= p12_data_enable ? p11_uge_4223 : p12_uge_4223;
      p12_uge_4298 <= p12_data_enable ? p11_uge_4298 : p12_uge_4298;
      p12_uge_4364 <= p12_data_enable ? p11_uge_4364 : p12_uge_4364;
      p12_uge_4430 <= p12_data_enable ? p11_uge_4430 : p12_uge_4430;
      p12_uge_4496 <= p12_data_enable ? p11_uge_4496 : p12_uge_4496;
      p12_uge_4562 <= p12_data_enable ? p11_uge_4562 : p12_uge_4562;
      p12_uge_4628 <= p12_data_enable ? p11_uge_4628 : p12_uge_4628;
      p12_uge_4694 <= p12_data_enable ? p11_uge_4694 : p12_uge_4694;
      p12_uge_4760 <= p12_data_enable ? p11_uge_4760 : p12_uge_4760;
      p12_concat_4825 <= p12_data_enable ? concat_4825 : p12_concat_4825;
      p12_uge_4826 <= p12_data_enable ? uge_4826 : p12_uge_4826;
      p12_bit_slice_4007 <= p12_data_enable ? p11_bit_slice_4007 : p12_bit_slice_4007;
      p12_bit_slice_4008 <= p12_data_enable ? p11_bit_slice_4008 : p12_bit_slice_4008;
      p12_bit_slice_4009 <= p12_data_enable ? p11_bit_slice_4009 : p12_bit_slice_4009;
      p12_bit_slice_4010 <= p12_data_enable ? p11_bit_slice_4010 : p12_bit_slice_4010;
      p12_bit_slice_4011 <= p12_data_enable ? p11_bit_slice_4011 : p12_bit_slice_4011;
      p12_bit_slice_4012 <= p12_data_enable ? p11_bit_slice_4012 : p12_bit_slice_4012;
      p12_bit_slice_4013 <= p12_data_enable ? p11_bit_slice_4013 : p12_bit_slice_4013;
      p12_bit_slice_4014 <= p12_data_enable ? p11_bit_slice_4014 : p12_bit_slice_4014;
      p12_bit_slice_4015 <= p12_data_enable ? p11_bit_slice_4015 : p12_bit_slice_4015;
      p12_bit_slice_4017 <= p12_data_enable ? p11_bit_slice_4017 : p12_bit_slice_4017;
      p12_bit_slice_4018 <= p12_data_enable ? p11_bit_slice_4018 : p12_bit_slice_4018;
      p12_flag_zero <= p12_data_enable ? p11_flag_zero : p12_flag_zero;
      p12_result_sign <= p12_data_enable ? p11_result_sign : p12_result_sign;
      p12_result_exp <= p12_data_enable ? p11_result_exp : p12_result_exp;
      p13_b_fraction <= p13_data_enable ? p12_b_fraction : p13_b_fraction;
      p13_uge_4144 <= p13_data_enable ? p12_uge_4144 : p13_uge_4144;
      p13_b_fractionivisor__1 <= p13_data_enable ? p12_b_fractionivisor__1 : p13_b_fractionivisor__1;
      p13_uge_4152 <= p13_data_enable ? p12_uge_4152 : p13_uge_4152;
      p13_uge_4223 <= p13_data_enable ? p12_uge_4223 : p13_uge_4223;
      p13_uge_4298 <= p13_data_enable ? p12_uge_4298 : p13_uge_4298;
      p13_uge_4364 <= p13_data_enable ? p12_uge_4364 : p13_uge_4364;
      p13_uge_4430 <= p13_data_enable ? p12_uge_4430 : p13_uge_4430;
      p13_uge_4496 <= p13_data_enable ? p12_uge_4496 : p13_uge_4496;
      p13_uge_4562 <= p13_data_enable ? p12_uge_4562 : p13_uge_4562;
      p13_uge_4628 <= p13_data_enable ? p12_uge_4628 : p13_uge_4628;
      p13_uge_4694 <= p13_data_enable ? p12_uge_4694 : p13_uge_4694;
      p13_uge_4760 <= p13_data_enable ? p12_uge_4760 : p13_uge_4760;
      p13_uge_4826 <= p13_data_enable ? p12_uge_4826 : p13_uge_4826;
      p13_concat_4891 <= p13_data_enable ? concat_4891 : p13_concat_4891;
      p13_uge_4892 <= p13_data_enable ? uge_4892 : p13_uge_4892;
      p13_bit_slice_4008 <= p13_data_enable ? p12_bit_slice_4008 : p13_bit_slice_4008;
      p13_bit_slice_4009 <= p13_data_enable ? p12_bit_slice_4009 : p13_bit_slice_4009;
      p13_bit_slice_4010 <= p13_data_enable ? p12_bit_slice_4010 : p13_bit_slice_4010;
      p13_bit_slice_4011 <= p13_data_enable ? p12_bit_slice_4011 : p13_bit_slice_4011;
      p13_bit_slice_4012 <= p13_data_enable ? p12_bit_slice_4012 : p13_bit_slice_4012;
      p13_bit_slice_4013 <= p13_data_enable ? p12_bit_slice_4013 : p13_bit_slice_4013;
      p13_bit_slice_4014 <= p13_data_enable ? p12_bit_slice_4014 : p13_bit_slice_4014;
      p13_bit_slice_4015 <= p13_data_enable ? p12_bit_slice_4015 : p13_bit_slice_4015;
      p13_bit_slice_4017 <= p13_data_enable ? p12_bit_slice_4017 : p13_bit_slice_4017;
      p13_bit_slice_4018 <= p13_data_enable ? p12_bit_slice_4018 : p13_bit_slice_4018;
      p13_flag_zero <= p13_data_enable ? p12_flag_zero : p13_flag_zero;
      p13_result_sign <= p13_data_enable ? p12_result_sign : p13_result_sign;
      p13_result_exp <= p13_data_enable ? p12_result_exp : p13_result_exp;
      p14_b_fraction <= p14_data_enable ? p13_b_fraction : p14_b_fraction;
      p14_uge_4144 <= p14_data_enable ? p13_uge_4144 : p14_uge_4144;
      p14_b_fractionivisor__1 <= p14_data_enable ? p13_b_fractionivisor__1 : p14_b_fractionivisor__1;
      p14_uge_4152 <= p14_data_enable ? p13_uge_4152 : p14_uge_4152;
      p14_uge_4223 <= p14_data_enable ? p13_uge_4223 : p14_uge_4223;
      p14_uge_4298 <= p14_data_enable ? p13_uge_4298 : p14_uge_4298;
      p14_uge_4364 <= p14_data_enable ? p13_uge_4364 : p14_uge_4364;
      p14_uge_4430 <= p14_data_enable ? p13_uge_4430 : p14_uge_4430;
      p14_uge_4496 <= p14_data_enable ? p13_uge_4496 : p14_uge_4496;
      p14_uge_4562 <= p14_data_enable ? p13_uge_4562 : p14_uge_4562;
      p14_uge_4628 <= p14_data_enable ? p13_uge_4628 : p14_uge_4628;
      p14_uge_4694 <= p14_data_enable ? p13_uge_4694 : p14_uge_4694;
      p14_uge_4760 <= p14_data_enable ? p13_uge_4760 : p14_uge_4760;
      p14_uge_4826 <= p14_data_enable ? p13_uge_4826 : p14_uge_4826;
      p14_uge_4892 <= p14_data_enable ? p13_uge_4892 : p14_uge_4892;
      p14_concat_4957 <= p14_data_enable ? concat_4957 : p14_concat_4957;
      p14_uge_4958 <= p14_data_enable ? uge_4958 : p14_uge_4958;
      p14_bit_slice_4009 <= p14_data_enable ? p13_bit_slice_4009 : p14_bit_slice_4009;
      p14_bit_slice_4010 <= p14_data_enable ? p13_bit_slice_4010 : p14_bit_slice_4010;
      p14_bit_slice_4011 <= p14_data_enable ? p13_bit_slice_4011 : p14_bit_slice_4011;
      p14_bit_slice_4012 <= p14_data_enable ? p13_bit_slice_4012 : p14_bit_slice_4012;
      p14_bit_slice_4013 <= p14_data_enable ? p13_bit_slice_4013 : p14_bit_slice_4013;
      p14_bit_slice_4014 <= p14_data_enable ? p13_bit_slice_4014 : p14_bit_slice_4014;
      p14_bit_slice_4015 <= p14_data_enable ? p13_bit_slice_4015 : p14_bit_slice_4015;
      p14_bit_slice_4017 <= p14_data_enable ? p13_bit_slice_4017 : p14_bit_slice_4017;
      p14_bit_slice_4018 <= p14_data_enable ? p13_bit_slice_4018 : p14_bit_slice_4018;
      p14_flag_zero <= p14_data_enable ? p13_flag_zero : p14_flag_zero;
      p14_result_sign <= p14_data_enable ? p13_result_sign : p14_result_sign;
      p14_result_exp <= p14_data_enable ? p13_result_exp : p14_result_exp;
      p15_b_fraction <= p15_data_enable ? p14_b_fraction : p15_b_fraction;
      p15_uge_4144 <= p15_data_enable ? p14_uge_4144 : p15_uge_4144;
      p15_b_fractionivisor__1 <= p15_data_enable ? p14_b_fractionivisor__1 : p15_b_fractionivisor__1;
      p15_uge_4152 <= p15_data_enable ? p14_uge_4152 : p15_uge_4152;
      p15_uge_4223 <= p15_data_enable ? p14_uge_4223 : p15_uge_4223;
      p15_uge_4298 <= p15_data_enable ? p14_uge_4298 : p15_uge_4298;
      p15_uge_4364 <= p15_data_enable ? p14_uge_4364 : p15_uge_4364;
      p15_uge_4430 <= p15_data_enable ? p14_uge_4430 : p15_uge_4430;
      p15_uge_4496 <= p15_data_enable ? p14_uge_4496 : p15_uge_4496;
      p15_uge_4562 <= p15_data_enable ? p14_uge_4562 : p15_uge_4562;
      p15_uge_4628 <= p15_data_enable ? p14_uge_4628 : p15_uge_4628;
      p15_uge_4694 <= p15_data_enable ? p14_uge_4694 : p15_uge_4694;
      p15_uge_4760 <= p15_data_enable ? p14_uge_4760 : p15_uge_4760;
      p15_uge_4826 <= p15_data_enable ? p14_uge_4826 : p15_uge_4826;
      p15_uge_4892 <= p15_data_enable ? p14_uge_4892 : p15_uge_4892;
      p15_uge_4958 <= p15_data_enable ? p14_uge_4958 : p15_uge_4958;
      p15_concat_5023 <= p15_data_enable ? concat_5023 : p15_concat_5023;
      p15_uge_5024 <= p15_data_enable ? uge_5024 : p15_uge_5024;
      p15_bit_slice_4010 <= p15_data_enable ? p14_bit_slice_4010 : p15_bit_slice_4010;
      p15_bit_slice_4011 <= p15_data_enable ? p14_bit_slice_4011 : p15_bit_slice_4011;
      p15_bit_slice_4012 <= p15_data_enable ? p14_bit_slice_4012 : p15_bit_slice_4012;
      p15_bit_slice_4013 <= p15_data_enable ? p14_bit_slice_4013 : p15_bit_slice_4013;
      p15_bit_slice_4014 <= p15_data_enable ? p14_bit_slice_4014 : p15_bit_slice_4014;
      p15_bit_slice_4015 <= p15_data_enable ? p14_bit_slice_4015 : p15_bit_slice_4015;
      p15_bit_slice_4017 <= p15_data_enable ? p14_bit_slice_4017 : p15_bit_slice_4017;
      p15_bit_slice_4018 <= p15_data_enable ? p14_bit_slice_4018 : p15_bit_slice_4018;
      p15_flag_zero <= p15_data_enable ? p14_flag_zero : p15_flag_zero;
      p15_result_sign <= p15_data_enable ? p14_result_sign : p15_result_sign;
      p15_result_exp <= p15_data_enable ? p14_result_exp : p15_result_exp;
      p16_b_fraction <= p16_data_enable ? p15_b_fraction : p16_b_fraction;
      p16_uge_4144 <= p16_data_enable ? p15_uge_4144 : p16_uge_4144;
      p16_b_fractionivisor__1 <= p16_data_enable ? p15_b_fractionivisor__1 : p16_b_fractionivisor__1;
      p16_uge_4152 <= p16_data_enable ? p15_uge_4152 : p16_uge_4152;
      p16_uge_4223 <= p16_data_enable ? p15_uge_4223 : p16_uge_4223;
      p16_uge_4298 <= p16_data_enable ? p15_uge_4298 : p16_uge_4298;
      p16_uge_4364 <= p16_data_enable ? p15_uge_4364 : p16_uge_4364;
      p16_uge_4430 <= p16_data_enable ? p15_uge_4430 : p16_uge_4430;
      p16_uge_4496 <= p16_data_enable ? p15_uge_4496 : p16_uge_4496;
      p16_uge_4562 <= p16_data_enable ? p15_uge_4562 : p16_uge_4562;
      p16_uge_4628 <= p16_data_enable ? p15_uge_4628 : p16_uge_4628;
      p16_uge_4694 <= p16_data_enable ? p15_uge_4694 : p16_uge_4694;
      p16_uge_4760 <= p16_data_enable ? p15_uge_4760 : p16_uge_4760;
      p16_uge_4826 <= p16_data_enable ? p15_uge_4826 : p16_uge_4826;
      p16_uge_4892 <= p16_data_enable ? p15_uge_4892 : p16_uge_4892;
      p16_uge_4958 <= p16_data_enable ? p15_uge_4958 : p16_uge_4958;
      p16_uge_5024 <= p16_data_enable ? p15_uge_5024 : p16_uge_5024;
      p16_concat_5089 <= p16_data_enable ? concat_5089 : p16_concat_5089;
      p16_uge_5090 <= p16_data_enable ? uge_5090 : p16_uge_5090;
      p16_bit_slice_4011 <= p16_data_enable ? p15_bit_slice_4011 : p16_bit_slice_4011;
      p16_bit_slice_4012 <= p16_data_enable ? p15_bit_slice_4012 : p16_bit_slice_4012;
      p16_bit_slice_4013 <= p16_data_enable ? p15_bit_slice_4013 : p16_bit_slice_4013;
      p16_bit_slice_4014 <= p16_data_enable ? p15_bit_slice_4014 : p16_bit_slice_4014;
      p16_bit_slice_4015 <= p16_data_enable ? p15_bit_slice_4015 : p16_bit_slice_4015;
      p16_bit_slice_4017 <= p16_data_enable ? p15_bit_slice_4017 : p16_bit_slice_4017;
      p16_bit_slice_4018 <= p16_data_enable ? p15_bit_slice_4018 : p16_bit_slice_4018;
      p16_flag_zero <= p16_data_enable ? p15_flag_zero : p16_flag_zero;
      p16_result_sign <= p16_data_enable ? p15_result_sign : p16_result_sign;
      p16_result_exp <= p16_data_enable ? p15_result_exp : p16_result_exp;
      p17_b_fraction <= p17_data_enable ? p16_b_fraction : p17_b_fraction;
      p17_uge_4144 <= p17_data_enable ? p16_uge_4144 : p17_uge_4144;
      p17_b_fractionivisor__1 <= p17_data_enable ? p16_b_fractionivisor__1 : p17_b_fractionivisor__1;
      p17_uge_4152 <= p17_data_enable ? p16_uge_4152 : p17_uge_4152;
      p17_uge_4223 <= p17_data_enable ? p16_uge_4223 : p17_uge_4223;
      p17_uge_4298 <= p17_data_enable ? p16_uge_4298 : p17_uge_4298;
      p17_uge_4364 <= p17_data_enable ? p16_uge_4364 : p17_uge_4364;
      p17_uge_4430 <= p17_data_enable ? p16_uge_4430 : p17_uge_4430;
      p17_uge_4496 <= p17_data_enable ? p16_uge_4496 : p17_uge_4496;
      p17_uge_4562 <= p17_data_enable ? p16_uge_4562 : p17_uge_4562;
      p17_uge_4628 <= p17_data_enable ? p16_uge_4628 : p17_uge_4628;
      p17_uge_4694 <= p17_data_enable ? p16_uge_4694 : p17_uge_4694;
      p17_uge_4760 <= p17_data_enable ? p16_uge_4760 : p17_uge_4760;
      p17_uge_4826 <= p17_data_enable ? p16_uge_4826 : p17_uge_4826;
      p17_uge_4892 <= p17_data_enable ? p16_uge_4892 : p17_uge_4892;
      p17_uge_4958 <= p17_data_enable ? p16_uge_4958 : p17_uge_4958;
      p17_uge_5024 <= p17_data_enable ? p16_uge_5024 : p17_uge_5024;
      p17_uge_5090 <= p17_data_enable ? p16_uge_5090 : p17_uge_5090;
      p17_concat_5155 <= p17_data_enable ? concat_5155 : p17_concat_5155;
      p17_uge_5156 <= p17_data_enable ? uge_5156 : p17_uge_5156;
      p17_bit_slice_4012 <= p17_data_enable ? p16_bit_slice_4012 : p17_bit_slice_4012;
      p17_bit_slice_4013 <= p17_data_enable ? p16_bit_slice_4013 : p17_bit_slice_4013;
      p17_bit_slice_4014 <= p17_data_enable ? p16_bit_slice_4014 : p17_bit_slice_4014;
      p17_bit_slice_4015 <= p17_data_enable ? p16_bit_slice_4015 : p17_bit_slice_4015;
      p17_bit_slice_4017 <= p17_data_enable ? p16_bit_slice_4017 : p17_bit_slice_4017;
      p17_bit_slice_4018 <= p17_data_enable ? p16_bit_slice_4018 : p17_bit_slice_4018;
      p17_flag_zero <= p17_data_enable ? p16_flag_zero : p17_flag_zero;
      p17_result_sign <= p17_data_enable ? p16_result_sign : p17_result_sign;
      p17_result_exp <= p17_data_enable ? p16_result_exp : p17_result_exp;
      p18_b_fraction <= p18_data_enable ? p17_b_fraction : p18_b_fraction;
      p18_uge_4144 <= p18_data_enable ? p17_uge_4144 : p18_uge_4144;
      p18_b_fractionivisor__1 <= p18_data_enable ? p17_b_fractionivisor__1 : p18_b_fractionivisor__1;
      p18_uge_4152 <= p18_data_enable ? p17_uge_4152 : p18_uge_4152;
      p18_uge_4223 <= p18_data_enable ? p17_uge_4223 : p18_uge_4223;
      p18_uge_4298 <= p18_data_enable ? p17_uge_4298 : p18_uge_4298;
      p18_uge_4364 <= p18_data_enable ? p17_uge_4364 : p18_uge_4364;
      p18_uge_4430 <= p18_data_enable ? p17_uge_4430 : p18_uge_4430;
      p18_uge_4496 <= p18_data_enable ? p17_uge_4496 : p18_uge_4496;
      p18_uge_4562 <= p18_data_enable ? p17_uge_4562 : p18_uge_4562;
      p18_uge_4628 <= p18_data_enable ? p17_uge_4628 : p18_uge_4628;
      p18_uge_4694 <= p18_data_enable ? p17_uge_4694 : p18_uge_4694;
      p18_uge_4760 <= p18_data_enable ? p17_uge_4760 : p18_uge_4760;
      p18_uge_4826 <= p18_data_enable ? p17_uge_4826 : p18_uge_4826;
      p18_uge_4892 <= p18_data_enable ? p17_uge_4892 : p18_uge_4892;
      p18_uge_4958 <= p18_data_enable ? p17_uge_4958 : p18_uge_4958;
      p18_uge_5024 <= p18_data_enable ? p17_uge_5024 : p18_uge_5024;
      p18_uge_5090 <= p18_data_enable ? p17_uge_5090 : p18_uge_5090;
      p18_uge_5156 <= p18_data_enable ? p17_uge_5156 : p18_uge_5156;
      p18_concat_5221 <= p18_data_enable ? concat_5221 : p18_concat_5221;
      p18_uge_5222 <= p18_data_enable ? uge_5222 : p18_uge_5222;
      p18_bit_slice_4013 <= p18_data_enable ? p17_bit_slice_4013 : p18_bit_slice_4013;
      p18_bit_slice_4014 <= p18_data_enable ? p17_bit_slice_4014 : p18_bit_slice_4014;
      p18_bit_slice_4015 <= p18_data_enable ? p17_bit_slice_4015 : p18_bit_slice_4015;
      p18_bit_slice_4017 <= p18_data_enable ? p17_bit_slice_4017 : p18_bit_slice_4017;
      p18_bit_slice_4018 <= p18_data_enable ? p17_bit_slice_4018 : p18_bit_slice_4018;
      p18_flag_zero <= p18_data_enable ? p17_flag_zero : p18_flag_zero;
      p18_result_sign <= p18_data_enable ? p17_result_sign : p18_result_sign;
      p18_result_exp <= p18_data_enable ? p17_result_exp : p18_result_exp;
      p19_b_fraction <= p19_data_enable ? p18_b_fraction : p19_b_fraction;
      p19_uge_4144 <= p19_data_enable ? p18_uge_4144 : p19_uge_4144;
      p19_b_fractionivisor__1 <= p19_data_enable ? p18_b_fractionivisor__1 : p19_b_fractionivisor__1;
      p19_uge_4152 <= p19_data_enable ? p18_uge_4152 : p19_uge_4152;
      p19_uge_4223 <= p19_data_enable ? p18_uge_4223 : p19_uge_4223;
      p19_uge_4298 <= p19_data_enable ? p18_uge_4298 : p19_uge_4298;
      p19_uge_4364 <= p19_data_enable ? p18_uge_4364 : p19_uge_4364;
      p19_uge_4430 <= p19_data_enable ? p18_uge_4430 : p19_uge_4430;
      p19_uge_4496 <= p19_data_enable ? p18_uge_4496 : p19_uge_4496;
      p19_uge_4562 <= p19_data_enable ? p18_uge_4562 : p19_uge_4562;
      p19_uge_4628 <= p19_data_enable ? p18_uge_4628 : p19_uge_4628;
      p19_uge_4694 <= p19_data_enable ? p18_uge_4694 : p19_uge_4694;
      p19_uge_4760 <= p19_data_enable ? p18_uge_4760 : p19_uge_4760;
      p19_uge_4826 <= p19_data_enable ? p18_uge_4826 : p19_uge_4826;
      p19_uge_4892 <= p19_data_enable ? p18_uge_4892 : p19_uge_4892;
      p19_uge_4958 <= p19_data_enable ? p18_uge_4958 : p19_uge_4958;
      p19_uge_5024 <= p19_data_enable ? p18_uge_5024 : p19_uge_5024;
      p19_uge_5090 <= p19_data_enable ? p18_uge_5090 : p19_uge_5090;
      p19_uge_5156 <= p19_data_enable ? p18_uge_5156 : p19_uge_5156;
      p19_uge_5222 <= p19_data_enable ? p18_uge_5222 : p19_uge_5222;
      p19_concat_5287 <= p19_data_enable ? concat_5287 : p19_concat_5287;
      p19_uge_5288 <= p19_data_enable ? uge_5288 : p19_uge_5288;
      p19_bit_slice_4014 <= p19_data_enable ? p18_bit_slice_4014 : p19_bit_slice_4014;
      p19_bit_slice_4015 <= p19_data_enable ? p18_bit_slice_4015 : p19_bit_slice_4015;
      p19_bit_slice_4017 <= p19_data_enable ? p18_bit_slice_4017 : p19_bit_slice_4017;
      p19_bit_slice_4018 <= p19_data_enable ? p18_bit_slice_4018 : p19_bit_slice_4018;
      p19_flag_zero <= p19_data_enable ? p18_flag_zero : p19_flag_zero;
      p19_result_sign <= p19_data_enable ? p18_result_sign : p19_result_sign;
      p19_result_exp <= p19_data_enable ? p18_result_exp : p19_result_exp;
      p20_b_fraction <= p20_data_enable ? p19_b_fraction : p20_b_fraction;
      p20_uge_4144 <= p20_data_enable ? p19_uge_4144 : p20_uge_4144;
      p20_b_fractionivisor__1 <= p20_data_enable ? p19_b_fractionivisor__1 : p20_b_fractionivisor__1;
      p20_uge_4152 <= p20_data_enable ? p19_uge_4152 : p20_uge_4152;
      p20_uge_4223 <= p20_data_enable ? p19_uge_4223 : p20_uge_4223;
      p20_uge_4298 <= p20_data_enable ? p19_uge_4298 : p20_uge_4298;
      p20_uge_4364 <= p20_data_enable ? p19_uge_4364 : p20_uge_4364;
      p20_uge_4430 <= p20_data_enable ? p19_uge_4430 : p20_uge_4430;
      p20_uge_4496 <= p20_data_enable ? p19_uge_4496 : p20_uge_4496;
      p20_uge_4562 <= p20_data_enable ? p19_uge_4562 : p20_uge_4562;
      p20_uge_4628 <= p20_data_enable ? p19_uge_4628 : p20_uge_4628;
      p20_uge_4694 <= p20_data_enable ? p19_uge_4694 : p20_uge_4694;
      p20_uge_4760 <= p20_data_enable ? p19_uge_4760 : p20_uge_4760;
      p20_uge_4826 <= p20_data_enable ? p19_uge_4826 : p20_uge_4826;
      p20_uge_4892 <= p20_data_enable ? p19_uge_4892 : p20_uge_4892;
      p20_uge_4958 <= p20_data_enable ? p19_uge_4958 : p20_uge_4958;
      p20_uge_5024 <= p20_data_enable ? p19_uge_5024 : p20_uge_5024;
      p20_uge_5090 <= p20_data_enable ? p19_uge_5090 : p20_uge_5090;
      p20_uge_5156 <= p20_data_enable ? p19_uge_5156 : p20_uge_5156;
      p20_uge_5222 <= p20_data_enable ? p19_uge_5222 : p20_uge_5222;
      p20_uge_5288 <= p20_data_enable ? p19_uge_5288 : p20_uge_5288;
      p20_concat_5353 <= p20_data_enable ? concat_5353 : p20_concat_5353;
      p20_uge_5354 <= p20_data_enable ? uge_5354 : p20_uge_5354;
      p20_bit_slice_4015 <= p20_data_enable ? p19_bit_slice_4015 : p20_bit_slice_4015;
      p20_bit_slice_4017 <= p20_data_enable ? p19_bit_slice_4017 : p20_bit_slice_4017;
      p20_bit_slice_4018 <= p20_data_enable ? p19_bit_slice_4018 : p20_bit_slice_4018;
      p20_flag_zero <= p20_data_enable ? p19_flag_zero : p20_flag_zero;
      p20_result_sign <= p20_data_enable ? p19_result_sign : p20_result_sign;
      p20_result_exp <= p20_data_enable ? p19_result_exp : p20_result_exp;
      p21_b_fraction <= p21_data_enable ? p20_b_fraction : p21_b_fraction;
      p21_uge_4144 <= p21_data_enable ? p20_uge_4144 : p21_uge_4144;
      p21_b_fractionivisor__1 <= p21_data_enable ? p20_b_fractionivisor__1 : p21_b_fractionivisor__1;
      p21_uge_4152 <= p21_data_enable ? p20_uge_4152 : p21_uge_4152;
      p21_uge_4223 <= p21_data_enable ? p20_uge_4223 : p21_uge_4223;
      p21_uge_4298 <= p21_data_enable ? p20_uge_4298 : p21_uge_4298;
      p21_uge_4364 <= p21_data_enable ? p20_uge_4364 : p21_uge_4364;
      p21_uge_4430 <= p21_data_enable ? p20_uge_4430 : p21_uge_4430;
      p21_uge_4496 <= p21_data_enable ? p20_uge_4496 : p21_uge_4496;
      p21_uge_4562 <= p21_data_enable ? p20_uge_4562 : p21_uge_4562;
      p21_uge_4628 <= p21_data_enable ? p20_uge_4628 : p21_uge_4628;
      p21_uge_4694 <= p21_data_enable ? p20_uge_4694 : p21_uge_4694;
      p21_uge_4760 <= p21_data_enable ? p20_uge_4760 : p21_uge_4760;
      p21_uge_4826 <= p21_data_enable ? p20_uge_4826 : p21_uge_4826;
      p21_uge_4892 <= p21_data_enable ? p20_uge_4892 : p21_uge_4892;
      p21_uge_4958 <= p21_data_enable ? p20_uge_4958 : p21_uge_4958;
      p21_uge_5024 <= p21_data_enable ? p20_uge_5024 : p21_uge_5024;
      p21_uge_5090 <= p21_data_enable ? p20_uge_5090 : p21_uge_5090;
      p21_uge_5156 <= p21_data_enable ? p20_uge_5156 : p21_uge_5156;
      p21_uge_5222 <= p21_data_enable ? p20_uge_5222 : p21_uge_5222;
      p21_uge_5288 <= p21_data_enable ? p20_uge_5288 : p21_uge_5288;
      p21_uge_5354 <= p21_data_enable ? p20_uge_5354 : p21_uge_5354;
      p21_concat_5419 <= p21_data_enable ? concat_5419 : p21_concat_5419;
      p21_uge_5420 <= p21_data_enable ? uge_5420 : p21_uge_5420;
      p21_bit_slice_4017 <= p21_data_enable ? p20_bit_slice_4017 : p21_bit_slice_4017;
      p21_bit_slice_4018 <= p21_data_enable ? p20_bit_slice_4018 : p21_bit_slice_4018;
      p21_flag_zero <= p21_data_enable ? p20_flag_zero : p21_flag_zero;
      p21_result_sign <= p21_data_enable ? p20_result_sign : p21_result_sign;
      p21_result_exp <= p21_data_enable ? p20_result_exp : p21_result_exp;
      p22_b_fraction <= p22_data_enable ? p21_b_fraction : p22_b_fraction;
      p22_uge_4144 <= p22_data_enable ? p21_uge_4144 : p22_uge_4144;
      p22_b_fractionivisor__1 <= p22_data_enable ? p21_b_fractionivisor__1 : p22_b_fractionivisor__1;
      p22_uge_4152 <= p22_data_enable ? p21_uge_4152 : p22_uge_4152;
      p22_uge_4223 <= p22_data_enable ? p21_uge_4223 : p22_uge_4223;
      p22_uge_4298 <= p22_data_enable ? p21_uge_4298 : p22_uge_4298;
      p22_uge_4364 <= p22_data_enable ? p21_uge_4364 : p22_uge_4364;
      p22_uge_4430 <= p22_data_enable ? p21_uge_4430 : p22_uge_4430;
      p22_uge_4496 <= p22_data_enable ? p21_uge_4496 : p22_uge_4496;
      p22_uge_4562 <= p22_data_enable ? p21_uge_4562 : p22_uge_4562;
      p22_uge_4628 <= p22_data_enable ? p21_uge_4628 : p22_uge_4628;
      p22_uge_4694 <= p22_data_enable ? p21_uge_4694 : p22_uge_4694;
      p22_uge_4760 <= p22_data_enable ? p21_uge_4760 : p22_uge_4760;
      p22_uge_4826 <= p22_data_enable ? p21_uge_4826 : p22_uge_4826;
      p22_uge_4892 <= p22_data_enable ? p21_uge_4892 : p22_uge_4892;
      p22_uge_4958 <= p22_data_enable ? p21_uge_4958 : p22_uge_4958;
      p22_uge_5024 <= p22_data_enable ? p21_uge_5024 : p22_uge_5024;
      p22_uge_5090 <= p22_data_enable ? p21_uge_5090 : p22_uge_5090;
      p22_uge_5156 <= p22_data_enable ? p21_uge_5156 : p22_uge_5156;
      p22_uge_5222 <= p22_data_enable ? p21_uge_5222 : p22_uge_5222;
      p22_uge_5288 <= p22_data_enable ? p21_uge_5288 : p22_uge_5288;
      p22_uge_5354 <= p22_data_enable ? p21_uge_5354 : p22_uge_5354;
      p22_uge_5420 <= p22_data_enable ? p21_uge_5420 : p22_uge_5420;
      p22_concat_5485 <= p22_data_enable ? concat_5485 : p22_concat_5485;
      p22_uge_5486 <= p22_data_enable ? uge_5486 : p22_uge_5486;
      p22_bit_slice_4018 <= p22_data_enable ? p21_bit_slice_4018 : p22_bit_slice_4018;
      p22_flag_zero <= p22_data_enable ? p21_flag_zero : p22_flag_zero;
      p22_result_sign <= p22_data_enable ? p21_result_sign : p22_result_sign;
      p22_result_exp <= p22_data_enable ? p21_result_exp : p22_result_exp;
      p23_uge_4144 <= p23_data_enable ? p22_uge_4144 : p23_uge_4144;
      p23_uge_4152 <= p23_data_enable ? p22_uge_4152 : p23_uge_4152;
      p23_uge_4223 <= p23_data_enable ? p22_uge_4223 : p23_uge_4223;
      p23_uge_4298 <= p23_data_enable ? p22_uge_4298 : p23_uge_4298;
      p23_uge_4364 <= p23_data_enable ? p22_uge_4364 : p23_uge_4364;
      p23_uge_4430 <= p23_data_enable ? p22_uge_4430 : p23_uge_4430;
      p23_uge_4496 <= p23_data_enable ? p22_uge_4496 : p23_uge_4496;
      p23_uge_4562 <= p23_data_enable ? p22_uge_4562 : p23_uge_4562;
      p23_uge_4628 <= p23_data_enable ? p22_uge_4628 : p23_uge_4628;
      p23_uge_4694 <= p23_data_enable ? p22_uge_4694 : p23_uge_4694;
      p23_uge_4760 <= p23_data_enable ? p22_uge_4760 : p23_uge_4760;
      p23_uge_4826 <= p23_data_enable ? p22_uge_4826 : p23_uge_4826;
      p23_uge_4892 <= p23_data_enable ? p22_uge_4892 : p23_uge_4892;
      p23_uge_4958 <= p23_data_enable ? p22_uge_4958 : p23_uge_4958;
      p23_uge_5024 <= p23_data_enable ? p22_uge_5024 : p23_uge_5024;
      p23_uge_5090 <= p23_data_enable ? p22_uge_5090 : p23_uge_5090;
      p23_uge_5156 <= p23_data_enable ? p22_uge_5156 : p23_uge_5156;
      p23_uge_5222 <= p23_data_enable ? p22_uge_5222 : p23_uge_5222;
      p23_uge_5288 <= p23_data_enable ? p22_uge_5288 : p23_uge_5288;
      p23_uge_5354 <= p23_data_enable ? p22_uge_5354 : p23_uge_5354;
      p23_uge_5420 <= p23_data_enable ? p22_uge_5420 : p23_uge_5420;
      p23_uge_5486 <= p23_data_enable ? p22_uge_5486 : p23_uge_5486;
      p23_flag_zero <= p23_data_enable ? p22_flag_zero : p23_flag_zero;
      p23_q__23_squeezed_portion_0_width_1 <= p23_data_enable ? q__23_squeezed_portion_0_width_1 : p23_q__23_squeezed_portion_0_width_1;
      p23_result_sign <= p23_data_enable ? p22_result_sign : p23_result_sign;
      p23_result_exp <= p23_data_enable ? p22_result_exp : p23_result_exp;
      p0_valid <= p0_enable ? xls_float_ips__lhs_vld : p0_valid;
      p1_valid <= p1_enable ? p1_stage_done : p1_valid;
      p2_valid <= p2_enable ? p1_valid : p2_valid;
      p3_valid <= p3_enable ? p2_valid : p3_valid;
      p4_valid <= p4_enable ? p3_valid : p4_valid;
      p5_valid <= p5_enable ? p4_valid : p5_valid;
      p6_valid <= p6_enable ? p5_valid : p6_valid;
      p7_valid <= p7_enable ? p6_valid : p7_valid;
      p8_valid <= p8_enable ? p7_valid : p8_valid;
      p9_valid <= p9_enable ? p8_valid : p9_valid;
      p10_valid <= p10_enable ? p9_valid : p10_valid;
      p11_valid <= p11_enable ? p10_valid : p11_valid;
      p12_valid <= p12_enable ? p11_valid : p12_valid;
      p13_valid <= p13_enable ? p12_valid : p13_valid;
      p14_valid <= p14_enable ? p13_valid : p14_valid;
      p15_valid <= p15_enable ? p14_valid : p15_valid;
      p16_valid <= p16_enable ? p15_valid : p16_valid;
      p17_valid <= p17_enable ? p16_valid : p17_valid;
      p18_valid <= p18_enable ? p17_valid : p18_valid;
      p19_valid <= p19_enable ? p18_valid : p19_valid;
      p20_valid <= p20_enable ? p19_valid : p20_valid;
      p21_valid <= p21_enable ? p20_valid : p21_valid;
      p22_valid <= p22_enable ? p21_valid : p22_valid;
      p23_valid <= p23_enable ? p22_valid : p23_valid;
      p24_valid <= p24_enable ? p24_stage_done : p24_valid;
      p25_valid <= p25_enable ? p24_valid : p25_valid;
      p26_valid <= p26_enable ? p25_valid : p26_valid;
      p27_valid <= p27_enable ? p26_valid : p27_valid;
      p28_valid <= p28_enable ? p27_valid : p28_valid;
      __xls_float_ips__result_reg <= xls_float_ips__result_load_en ? __xls_float_ips__result_buf : __xls_float_ips__result_reg;
      __xls_float_ips__result_valid_reg <= xls_float_ips__result_valid_load_en ? p23_valid : __xls_float_ips__result_valid_reg;
    end
  end
  assign xls_float_ips__result = __xls_float_ips__result_reg;
  assign xls_float_ips__result_vld = __xls_float_ips__result_valid_reg;
  assign xls_float_ips__lhs_rdy = p0_data_enable;
  assign xls_float_ips__rhs_rdy = p1_data_enable;
endmodule
module __xls_float_ips__divsi32_0_next(
  input wire clk,
  input wire rst,
  input wire [31:0] xls_float_ips__lhs,
  input wire xls_float_ips__lhs_vld,
  input wire [31:0] xls_float_ips__rhs,
  input wire xls_float_ips__rhs_vld,
  input wire xls_float_ips__result_rdy,
  output wire [31:0] xls_float_ips__result,
  output wire xls_float_ips__result_vld,
  output wire xls_float_ips__lhs_rdy,
  output wire xls_float_ips__rhs_rdy
);
  reg [31:0] p0_concat_6575;
  reg [31:0] p0_b;
  reg p0_bit_slice_6577;
  reg p0_bit_slice_6578;
  reg p0_bit_slice_6579;
  reg p0_bit_slice_6580;
  reg p0_bit_slice_6581;
  reg p0_bit_slice_6582;
  reg p0_bit_slice_6583;
  reg p0_bit_slice_6584;
  reg p0_bit_slice_6585;
  reg p0_bit_slice_6586;
  reg p0_bit_slice_6587;
  reg p0_bit_slice_6588;
  reg p0_bit_slice_6589;
  reg p0_bit_slice_6590;
  reg p0_bit_slice_6591;
  reg p0_bit_slice_6592;
  reg p0_bit_slice_6593;
  reg p0_bit_slice_6594;
  reg p0_bit_slice_6595;
  reg p0_bit_slice_6596;
  reg p0_bit_slice_6597;
  reg p0_bit_slice_6598;
  reg p0_bit_slice_6599;
  reg p0_bit_slice_6600;
  reg p0_bit_slice_6601;
  reg p0_bit_slice_6602;
  reg p0_bit_slice_6603;
  reg p0_bit_slice_6604;
  reg p0_bit_slice_6605;
  reg p0_bit_slice_6606;
  reg p0_bit_slice_6607;
  reg p0_negated;
  reg [31:0] p1_b;
  reg p1_uge_6683;
  reg [32:0] p1_bivisor__1;
  reg [31:0] p1_concat_6690;
  reg p1_uge_6691;
  reg p1_bit_slice_6578;
  reg p1_bit_slice_6579;
  reg p1_bit_slice_6580;
  reg p1_bit_slice_6581;
  reg p1_bit_slice_6582;
  reg p1_bit_slice_6583;
  reg p1_bit_slice_6584;
  reg p1_bit_slice_6585;
  reg p1_bit_slice_6586;
  reg p1_bit_slice_6587;
  reg p1_bit_slice_6588;
  reg p1_bit_slice_6589;
  reg p1_bit_slice_6590;
  reg p1_bit_slice_6591;
  reg p1_bit_slice_6592;
  reg p1_bit_slice_6593;
  reg p1_bit_slice_6594;
  reg p1_bit_slice_6595;
  reg p1_bit_slice_6596;
  reg p1_bit_slice_6597;
  reg p1_bit_slice_6598;
  reg p1_bit_slice_6599;
  reg p1_bit_slice_6600;
  reg p1_bit_slice_6601;
  reg p1_bit_slice_6602;
  reg p1_bit_slice_6603;
  reg p1_bit_slice_6604;
  reg p1_bit_slice_6605;
  reg p1_bit_slice_6606;
  reg p1_bit_slice_6607;
  reg p1_negated;
  reg [31:0] p2_b;
  reg p2_uge_6683;
  reg [32:0] p2_bivisor__1;
  reg p2_uge_6691;
  reg [31:0] p2_concat_6770;
  reg p2_uge_6771;
  reg p2_bit_slice_6579;
  reg p2_bit_slice_6580;
  reg p2_bit_slice_6581;
  reg p2_bit_slice_6582;
  reg p2_bit_slice_6583;
  reg p2_bit_slice_6584;
  reg p2_bit_slice_6585;
  reg p2_bit_slice_6586;
  reg p2_bit_slice_6587;
  reg p2_bit_slice_6588;
  reg p2_bit_slice_6589;
  reg p2_bit_slice_6590;
  reg p2_bit_slice_6591;
  reg p2_bit_slice_6592;
  reg p2_bit_slice_6593;
  reg p2_bit_slice_6594;
  reg p2_bit_slice_6595;
  reg p2_bit_slice_6596;
  reg p2_bit_slice_6597;
  reg p2_bit_slice_6598;
  reg p2_bit_slice_6599;
  reg p2_bit_slice_6600;
  reg p2_bit_slice_6601;
  reg p2_bit_slice_6602;
  reg p2_bit_slice_6603;
  reg p2_bit_slice_6604;
  reg p2_bit_slice_6605;
  reg p2_bit_slice_6606;
  reg p2_bit_slice_6607;
  reg p2_negated;
  reg [31:0] p3_b;
  reg p3_uge_6683;
  reg [32:0] p3_bivisor__1;
  reg p3_uge_6691;
  reg p3_uge_6771;
  reg [31:0] p3_concat_6850;
  reg p3_uge_6851;
  reg p3_bit_slice_6580;
  reg p3_bit_slice_6581;
  reg p3_bit_slice_6582;
  reg p3_bit_slice_6583;
  reg p3_bit_slice_6584;
  reg p3_bit_slice_6585;
  reg p3_bit_slice_6586;
  reg p3_bit_slice_6587;
  reg p3_bit_slice_6588;
  reg p3_bit_slice_6589;
  reg p3_bit_slice_6590;
  reg p3_bit_slice_6591;
  reg p3_bit_slice_6592;
  reg p3_bit_slice_6593;
  reg p3_bit_slice_6594;
  reg p3_bit_slice_6595;
  reg p3_bit_slice_6596;
  reg p3_bit_slice_6597;
  reg p3_bit_slice_6598;
  reg p3_bit_slice_6599;
  reg p3_bit_slice_6600;
  reg p3_bit_slice_6601;
  reg p3_bit_slice_6602;
  reg p3_bit_slice_6603;
  reg p3_bit_slice_6604;
  reg p3_bit_slice_6605;
  reg p3_bit_slice_6606;
  reg p3_bit_slice_6607;
  reg p3_negated;
  reg [31:0] p4_b;
  reg p4_uge_6683;
  reg [32:0] p4_bivisor__1;
  reg p4_uge_6691;
  reg p4_uge_6771;
  reg p4_uge_6851;
  reg [31:0] p4_concat_6930;
  reg p4_uge_6931;
  reg p4_bit_slice_6581;
  reg p4_bit_slice_6582;
  reg p4_bit_slice_6583;
  reg p4_bit_slice_6584;
  reg p4_bit_slice_6585;
  reg p4_bit_slice_6586;
  reg p4_bit_slice_6587;
  reg p4_bit_slice_6588;
  reg p4_bit_slice_6589;
  reg p4_bit_slice_6590;
  reg p4_bit_slice_6591;
  reg p4_bit_slice_6592;
  reg p4_bit_slice_6593;
  reg p4_bit_slice_6594;
  reg p4_bit_slice_6595;
  reg p4_bit_slice_6596;
  reg p4_bit_slice_6597;
  reg p4_bit_slice_6598;
  reg p4_bit_slice_6599;
  reg p4_bit_slice_6600;
  reg p4_bit_slice_6601;
  reg p4_bit_slice_6602;
  reg p4_bit_slice_6603;
  reg p4_bit_slice_6604;
  reg p4_bit_slice_6605;
  reg p4_bit_slice_6606;
  reg p4_bit_slice_6607;
  reg p4_negated;
  reg [31:0] p5_b;
  reg p5_uge_6683;
  reg [32:0] p5_bivisor__1;
  reg p5_uge_6691;
  reg p5_uge_6771;
  reg p5_uge_6851;
  reg p5_uge_6931;
  reg [31:0] p5_concat_7010;
  reg p5_uge_7011;
  reg p5_bit_slice_6582;
  reg p5_bit_slice_6583;
  reg p5_bit_slice_6584;
  reg p5_bit_slice_6585;
  reg p5_bit_slice_6586;
  reg p5_bit_slice_6587;
  reg p5_bit_slice_6588;
  reg p5_bit_slice_6589;
  reg p5_bit_slice_6590;
  reg p5_bit_slice_6591;
  reg p5_bit_slice_6592;
  reg p5_bit_slice_6593;
  reg p5_bit_slice_6594;
  reg p5_bit_slice_6595;
  reg p5_bit_slice_6596;
  reg p5_bit_slice_6597;
  reg p5_bit_slice_6598;
  reg p5_bit_slice_6599;
  reg p5_bit_slice_6600;
  reg p5_bit_slice_6601;
  reg p5_bit_slice_6602;
  reg p5_bit_slice_6603;
  reg p5_bit_slice_6604;
  reg p5_bit_slice_6605;
  reg p5_bit_slice_6606;
  reg p5_bit_slice_6607;
  reg p5_negated;
  reg [31:0] p6_b;
  reg p6_uge_6683;
  reg [32:0] p6_bivisor__1;
  reg p6_uge_6691;
  reg p6_uge_6771;
  reg p6_uge_6851;
  reg p6_uge_6931;
  reg p6_uge_7011;
  reg [31:0] p6_concat_7090;
  reg p6_uge_7091;
  reg p6_bit_slice_6583;
  reg p6_bit_slice_6584;
  reg p6_bit_slice_6585;
  reg p6_bit_slice_6586;
  reg p6_bit_slice_6587;
  reg p6_bit_slice_6588;
  reg p6_bit_slice_6589;
  reg p6_bit_slice_6590;
  reg p6_bit_slice_6591;
  reg p6_bit_slice_6592;
  reg p6_bit_slice_6593;
  reg p6_bit_slice_6594;
  reg p6_bit_slice_6595;
  reg p6_bit_slice_6596;
  reg p6_bit_slice_6597;
  reg p6_bit_slice_6598;
  reg p6_bit_slice_6599;
  reg p6_bit_slice_6600;
  reg p6_bit_slice_6601;
  reg p6_bit_slice_6602;
  reg p6_bit_slice_6603;
  reg p6_bit_slice_6604;
  reg p6_bit_slice_6605;
  reg p6_bit_slice_6606;
  reg p6_bit_slice_6607;
  reg p6_negated;
  reg [31:0] p7_b;
  reg p7_uge_6683;
  reg [32:0] p7_bivisor__1;
  reg p7_uge_6691;
  reg p7_uge_6771;
  reg p7_uge_6851;
  reg p7_uge_6931;
  reg p7_uge_7011;
  reg p7_uge_7091;
  reg [31:0] p7_concat_7170;
  reg p7_uge_7171;
  reg p7_bit_slice_6584;
  reg p7_bit_slice_6585;
  reg p7_bit_slice_6586;
  reg p7_bit_slice_6587;
  reg p7_bit_slice_6588;
  reg p7_bit_slice_6589;
  reg p7_bit_slice_6590;
  reg p7_bit_slice_6591;
  reg p7_bit_slice_6592;
  reg p7_bit_slice_6593;
  reg p7_bit_slice_6594;
  reg p7_bit_slice_6595;
  reg p7_bit_slice_6596;
  reg p7_bit_slice_6597;
  reg p7_bit_slice_6598;
  reg p7_bit_slice_6599;
  reg p7_bit_slice_6600;
  reg p7_bit_slice_6601;
  reg p7_bit_slice_6602;
  reg p7_bit_slice_6603;
  reg p7_bit_slice_6604;
  reg p7_bit_slice_6605;
  reg p7_bit_slice_6606;
  reg p7_bit_slice_6607;
  reg p7_negated;
  reg [31:0] p8_b;
  reg p8_uge_6683;
  reg [32:0] p8_bivisor__1;
  reg p8_uge_6691;
  reg p8_uge_6771;
  reg p8_uge_6851;
  reg p8_uge_6931;
  reg p8_uge_7011;
  reg p8_uge_7091;
  reg p8_uge_7171;
  reg [31:0] p8_concat_7250;
  reg p8_uge_7251;
  reg p8_bit_slice_6585;
  reg p8_bit_slice_6586;
  reg p8_bit_slice_6587;
  reg p8_bit_slice_6588;
  reg p8_bit_slice_6589;
  reg p8_bit_slice_6590;
  reg p8_bit_slice_6591;
  reg p8_bit_slice_6592;
  reg p8_bit_slice_6593;
  reg p8_bit_slice_6594;
  reg p8_bit_slice_6595;
  reg p8_bit_slice_6596;
  reg p8_bit_slice_6597;
  reg p8_bit_slice_6598;
  reg p8_bit_slice_6599;
  reg p8_bit_slice_6600;
  reg p8_bit_slice_6601;
  reg p8_bit_slice_6602;
  reg p8_bit_slice_6603;
  reg p8_bit_slice_6604;
  reg p8_bit_slice_6605;
  reg p8_bit_slice_6606;
  reg p8_bit_slice_6607;
  reg p8_negated;
  reg [31:0] p9_b;
  reg p9_uge_6683;
  reg [32:0] p9_bivisor__1;
  reg p9_uge_6691;
  reg p9_uge_6771;
  reg p9_uge_6851;
  reg p9_uge_6931;
  reg p9_uge_7011;
  reg p9_uge_7091;
  reg p9_uge_7171;
  reg p9_uge_7251;
  reg [31:0] p9_concat_7330;
  reg p9_uge_7331;
  reg p9_bit_slice_6586;
  reg p9_bit_slice_6587;
  reg p9_bit_slice_6588;
  reg p9_bit_slice_6589;
  reg p9_bit_slice_6590;
  reg p9_bit_slice_6591;
  reg p9_bit_slice_6592;
  reg p9_bit_slice_6593;
  reg p9_bit_slice_6594;
  reg p9_bit_slice_6595;
  reg p9_bit_slice_6596;
  reg p9_bit_slice_6597;
  reg p9_bit_slice_6598;
  reg p9_bit_slice_6599;
  reg p9_bit_slice_6600;
  reg p9_bit_slice_6601;
  reg p9_bit_slice_6602;
  reg p9_bit_slice_6603;
  reg p9_bit_slice_6604;
  reg p9_bit_slice_6605;
  reg p9_bit_slice_6606;
  reg p9_bit_slice_6607;
  reg p9_negated;
  reg [31:0] p10_b;
  reg p10_uge_6683;
  reg [32:0] p10_bivisor__1;
  reg p10_uge_6691;
  reg p10_uge_6771;
  reg p10_uge_6851;
  reg p10_uge_6931;
  reg p10_uge_7011;
  reg p10_uge_7091;
  reg p10_uge_7171;
  reg p10_uge_7251;
  reg p10_uge_7331;
  reg [31:0] p10_concat_7410;
  reg p10_uge_7411;
  reg p10_bit_slice_6587;
  reg p10_bit_slice_6588;
  reg p10_bit_slice_6589;
  reg p10_bit_slice_6590;
  reg p10_bit_slice_6591;
  reg p10_bit_slice_6592;
  reg p10_bit_slice_6593;
  reg p10_bit_slice_6594;
  reg p10_bit_slice_6595;
  reg p10_bit_slice_6596;
  reg p10_bit_slice_6597;
  reg p10_bit_slice_6598;
  reg p10_bit_slice_6599;
  reg p10_bit_slice_6600;
  reg p10_bit_slice_6601;
  reg p10_bit_slice_6602;
  reg p10_bit_slice_6603;
  reg p10_bit_slice_6604;
  reg p10_bit_slice_6605;
  reg p10_bit_slice_6606;
  reg p10_bit_slice_6607;
  reg p10_negated;
  reg [31:0] p11_b;
  reg p11_uge_6683;
  reg [32:0] p11_bivisor__1;
  reg p11_uge_6691;
  reg p11_uge_6771;
  reg p11_uge_6851;
  reg p11_uge_6931;
  reg p11_uge_7011;
  reg p11_uge_7091;
  reg p11_uge_7171;
  reg p11_uge_7251;
  reg p11_uge_7331;
  reg p11_uge_7411;
  reg [31:0] p11_concat_7490;
  reg p11_uge_7491;
  reg p11_bit_slice_6588;
  reg p11_bit_slice_6589;
  reg p11_bit_slice_6590;
  reg p11_bit_slice_6591;
  reg p11_bit_slice_6592;
  reg p11_bit_slice_6593;
  reg p11_bit_slice_6594;
  reg p11_bit_slice_6595;
  reg p11_bit_slice_6596;
  reg p11_bit_slice_6597;
  reg p11_bit_slice_6598;
  reg p11_bit_slice_6599;
  reg p11_bit_slice_6600;
  reg p11_bit_slice_6601;
  reg p11_bit_slice_6602;
  reg p11_bit_slice_6603;
  reg p11_bit_slice_6604;
  reg p11_bit_slice_6605;
  reg p11_bit_slice_6606;
  reg p11_bit_slice_6607;
  reg p11_negated;
  reg [31:0] p12_b;
  reg p12_uge_6683;
  reg [32:0] p12_bivisor__1;
  reg p12_uge_6691;
  reg p12_uge_6771;
  reg p12_uge_6851;
  reg p12_uge_6931;
  reg p12_uge_7011;
  reg p12_uge_7091;
  reg p12_uge_7171;
  reg p12_uge_7251;
  reg p12_uge_7331;
  reg p12_uge_7411;
  reg p12_uge_7491;
  reg [31:0] p12_concat_7570;
  reg p12_uge_7571;
  reg p12_bit_slice_6589;
  reg p12_bit_slice_6590;
  reg p12_bit_slice_6591;
  reg p12_bit_slice_6592;
  reg p12_bit_slice_6593;
  reg p12_bit_slice_6594;
  reg p12_bit_slice_6595;
  reg p12_bit_slice_6596;
  reg p12_bit_slice_6597;
  reg p12_bit_slice_6598;
  reg p12_bit_slice_6599;
  reg p12_bit_slice_6600;
  reg p12_bit_slice_6601;
  reg p12_bit_slice_6602;
  reg p12_bit_slice_6603;
  reg p12_bit_slice_6604;
  reg p12_bit_slice_6605;
  reg p12_bit_slice_6606;
  reg p12_bit_slice_6607;
  reg p12_negated;
  reg [31:0] p13_b;
  reg p13_uge_6683;
  reg [32:0] p13_bivisor__1;
  reg p13_uge_6691;
  reg p13_uge_6771;
  reg p13_uge_6851;
  reg p13_uge_6931;
  reg p13_uge_7011;
  reg p13_uge_7091;
  reg p13_uge_7171;
  reg p13_uge_7251;
  reg p13_uge_7331;
  reg p13_uge_7411;
  reg p13_uge_7491;
  reg p13_uge_7571;
  reg [31:0] p13_concat_7650;
  reg p13_uge_7651;
  reg p13_bit_slice_6590;
  reg p13_bit_slice_6591;
  reg p13_bit_slice_6592;
  reg p13_bit_slice_6593;
  reg p13_bit_slice_6594;
  reg p13_bit_slice_6595;
  reg p13_bit_slice_6596;
  reg p13_bit_slice_6597;
  reg p13_bit_slice_6598;
  reg p13_bit_slice_6599;
  reg p13_bit_slice_6600;
  reg p13_bit_slice_6601;
  reg p13_bit_slice_6602;
  reg p13_bit_slice_6603;
  reg p13_bit_slice_6604;
  reg p13_bit_slice_6605;
  reg p13_bit_slice_6606;
  reg p13_bit_slice_6607;
  reg p13_negated;
  reg [31:0] p14_b;
  reg p14_uge_6683;
  reg [32:0] p14_bivisor__1;
  reg p14_uge_6691;
  reg p14_uge_6771;
  reg p14_uge_6851;
  reg p14_uge_6931;
  reg p14_uge_7011;
  reg p14_uge_7091;
  reg p14_uge_7171;
  reg p14_uge_7251;
  reg p14_uge_7331;
  reg p14_uge_7411;
  reg p14_uge_7491;
  reg p14_uge_7571;
  reg p14_uge_7651;
  reg [31:0] p14_concat_7730;
  reg p14_uge_7731;
  reg p14_bit_slice_6591;
  reg p14_bit_slice_6592;
  reg p14_bit_slice_6593;
  reg p14_bit_slice_6594;
  reg p14_bit_slice_6595;
  reg p14_bit_slice_6596;
  reg p14_bit_slice_6597;
  reg p14_bit_slice_6598;
  reg p14_bit_slice_6599;
  reg p14_bit_slice_6600;
  reg p14_bit_slice_6601;
  reg p14_bit_slice_6602;
  reg p14_bit_slice_6603;
  reg p14_bit_slice_6604;
  reg p14_bit_slice_6605;
  reg p14_bit_slice_6606;
  reg p14_bit_slice_6607;
  reg p14_negated;
  reg [31:0] p15_b;
  reg p15_uge_6683;
  reg [32:0] p15_bivisor__1;
  reg p15_uge_6691;
  reg p15_uge_6771;
  reg p15_uge_6851;
  reg p15_uge_6931;
  reg p15_uge_7011;
  reg p15_uge_7091;
  reg p15_uge_7171;
  reg p15_uge_7251;
  reg p15_uge_7331;
  reg p15_uge_7411;
  reg p15_uge_7491;
  reg p15_uge_7571;
  reg p15_uge_7651;
  reg p15_uge_7731;
  reg [31:0] p15_concat_7810;
  reg p15_uge_7811;
  reg p15_bit_slice_6592;
  reg p15_bit_slice_6593;
  reg p15_bit_slice_6594;
  reg p15_bit_slice_6595;
  reg p15_bit_slice_6596;
  reg p15_bit_slice_6597;
  reg p15_bit_slice_6598;
  reg p15_bit_slice_6599;
  reg p15_bit_slice_6600;
  reg p15_bit_slice_6601;
  reg p15_bit_slice_6602;
  reg p15_bit_slice_6603;
  reg p15_bit_slice_6604;
  reg p15_bit_slice_6605;
  reg p15_bit_slice_6606;
  reg p15_bit_slice_6607;
  reg p15_negated;
  reg [31:0] p16_b;
  reg p16_uge_6683;
  reg [32:0] p16_bivisor__1;
  reg p16_uge_6691;
  reg p16_uge_6771;
  reg p16_uge_6851;
  reg p16_uge_6931;
  reg p16_uge_7011;
  reg p16_uge_7091;
  reg p16_uge_7171;
  reg p16_uge_7251;
  reg p16_uge_7331;
  reg p16_uge_7411;
  reg p16_uge_7491;
  reg p16_uge_7571;
  reg p16_uge_7651;
  reg p16_uge_7731;
  reg p16_uge_7811;
  reg [31:0] p16_concat_7890;
  reg p16_uge_7891;
  reg p16_bit_slice_6593;
  reg p16_bit_slice_6594;
  reg p16_bit_slice_6595;
  reg p16_bit_slice_6596;
  reg p16_bit_slice_6597;
  reg p16_bit_slice_6598;
  reg p16_bit_slice_6599;
  reg p16_bit_slice_6600;
  reg p16_bit_slice_6601;
  reg p16_bit_slice_6602;
  reg p16_bit_slice_6603;
  reg p16_bit_slice_6604;
  reg p16_bit_slice_6605;
  reg p16_bit_slice_6606;
  reg p16_bit_slice_6607;
  reg p16_negated;
  reg [31:0] p17_b;
  reg p17_uge_6683;
  reg [32:0] p17_bivisor__1;
  reg p17_uge_6691;
  reg p17_uge_6771;
  reg p17_uge_6851;
  reg p17_uge_6931;
  reg p17_uge_7011;
  reg p17_uge_7091;
  reg p17_uge_7171;
  reg p17_uge_7251;
  reg p17_uge_7331;
  reg p17_uge_7411;
  reg p17_uge_7491;
  reg p17_uge_7571;
  reg p17_uge_7651;
  reg p17_uge_7731;
  reg p17_uge_7811;
  reg p17_uge_7891;
  reg [31:0] p17_concat_7970;
  reg p17_uge_7971;
  reg p17_bit_slice_6594;
  reg p17_bit_slice_6595;
  reg p17_bit_slice_6596;
  reg p17_bit_slice_6597;
  reg p17_bit_slice_6598;
  reg p17_bit_slice_6599;
  reg p17_bit_slice_6600;
  reg p17_bit_slice_6601;
  reg p17_bit_slice_6602;
  reg p17_bit_slice_6603;
  reg p17_bit_slice_6604;
  reg p17_bit_slice_6605;
  reg p17_bit_slice_6606;
  reg p17_bit_slice_6607;
  reg p17_negated;
  reg [31:0] p18_b;
  reg p18_uge_6683;
  reg [32:0] p18_bivisor__1;
  reg p18_uge_6691;
  reg p18_uge_6771;
  reg p18_uge_6851;
  reg p18_uge_6931;
  reg p18_uge_7011;
  reg p18_uge_7091;
  reg p18_uge_7171;
  reg p18_uge_7251;
  reg p18_uge_7331;
  reg p18_uge_7411;
  reg p18_uge_7491;
  reg p18_uge_7571;
  reg p18_uge_7651;
  reg p18_uge_7731;
  reg p18_uge_7811;
  reg p18_uge_7891;
  reg p18_uge_7971;
  reg [31:0] p18_concat_8050;
  reg p18_uge_8051;
  reg p18_bit_slice_6595;
  reg p18_bit_slice_6596;
  reg p18_bit_slice_6597;
  reg p18_bit_slice_6598;
  reg p18_bit_slice_6599;
  reg p18_bit_slice_6600;
  reg p18_bit_slice_6601;
  reg p18_bit_slice_6602;
  reg p18_bit_slice_6603;
  reg p18_bit_slice_6604;
  reg p18_bit_slice_6605;
  reg p18_bit_slice_6606;
  reg p18_bit_slice_6607;
  reg p18_negated;
  reg [31:0] p19_b;
  reg p19_uge_6683;
  reg [32:0] p19_bivisor__1;
  reg p19_uge_6691;
  reg p19_uge_6771;
  reg p19_uge_6851;
  reg p19_uge_6931;
  reg p19_uge_7011;
  reg p19_uge_7091;
  reg p19_uge_7171;
  reg p19_uge_7251;
  reg p19_uge_7331;
  reg p19_uge_7411;
  reg p19_uge_7491;
  reg p19_uge_7571;
  reg p19_uge_7651;
  reg p19_uge_7731;
  reg p19_uge_7811;
  reg p19_uge_7891;
  reg p19_uge_7971;
  reg p19_uge_8051;
  reg [31:0] p19_concat_8130;
  reg p19_uge_8131;
  reg p19_bit_slice_6596;
  reg p19_bit_slice_6597;
  reg p19_bit_slice_6598;
  reg p19_bit_slice_6599;
  reg p19_bit_slice_6600;
  reg p19_bit_slice_6601;
  reg p19_bit_slice_6602;
  reg p19_bit_slice_6603;
  reg p19_bit_slice_6604;
  reg p19_bit_slice_6605;
  reg p19_bit_slice_6606;
  reg p19_bit_slice_6607;
  reg p19_negated;
  reg [31:0] p20_b;
  reg p20_uge_6683;
  reg [32:0] p20_bivisor__1;
  reg p20_uge_6691;
  reg p20_uge_6771;
  reg p20_uge_6851;
  reg p20_uge_6931;
  reg p20_uge_7011;
  reg p20_uge_7091;
  reg p20_uge_7171;
  reg p20_uge_7251;
  reg p20_uge_7331;
  reg p20_uge_7411;
  reg p20_uge_7491;
  reg p20_uge_7571;
  reg p20_uge_7651;
  reg p20_uge_7731;
  reg p20_uge_7811;
  reg p20_uge_7891;
  reg p20_uge_7971;
  reg p20_uge_8051;
  reg p20_uge_8131;
  reg [31:0] p20_concat_8210;
  reg p20_uge_8211;
  reg p20_bit_slice_6597;
  reg p20_bit_slice_6598;
  reg p20_bit_slice_6599;
  reg p20_bit_slice_6600;
  reg p20_bit_slice_6601;
  reg p20_bit_slice_6602;
  reg p20_bit_slice_6603;
  reg p20_bit_slice_6604;
  reg p20_bit_slice_6605;
  reg p20_bit_slice_6606;
  reg p20_bit_slice_6607;
  reg p20_negated;
  reg [31:0] p21_b;
  reg p21_uge_6683;
  reg [32:0] p21_bivisor__1;
  reg p21_uge_6691;
  reg p21_uge_6771;
  reg p21_uge_6851;
  reg p21_uge_6931;
  reg p21_uge_7011;
  reg p21_uge_7091;
  reg p21_uge_7171;
  reg p21_uge_7251;
  reg p21_uge_7331;
  reg p21_uge_7411;
  reg p21_uge_7491;
  reg p21_uge_7571;
  reg p21_uge_7651;
  reg p21_uge_7731;
  reg p21_uge_7811;
  reg p21_uge_7891;
  reg p21_uge_7971;
  reg p21_uge_8051;
  reg p21_uge_8131;
  reg p21_uge_8211;
  reg [31:0] p21_concat_8290;
  reg p21_uge_8291;
  reg p21_bit_slice_6598;
  reg p21_bit_slice_6599;
  reg p21_bit_slice_6600;
  reg p21_bit_slice_6601;
  reg p21_bit_slice_6602;
  reg p21_bit_slice_6603;
  reg p21_bit_slice_6604;
  reg p21_bit_slice_6605;
  reg p21_bit_slice_6606;
  reg p21_bit_slice_6607;
  reg p21_negated;
  reg [31:0] p22_b;
  reg p22_uge_6683;
  reg [32:0] p22_bivisor__1;
  reg p22_uge_6691;
  reg p22_uge_6771;
  reg p22_uge_6851;
  reg p22_uge_6931;
  reg p22_uge_7011;
  reg p22_uge_7091;
  reg p22_uge_7171;
  reg p22_uge_7251;
  reg p22_uge_7331;
  reg p22_uge_7411;
  reg p22_uge_7491;
  reg p22_uge_7571;
  reg p22_uge_7651;
  reg p22_uge_7731;
  reg p22_uge_7811;
  reg p22_uge_7891;
  reg p22_uge_7971;
  reg p22_uge_8051;
  reg p22_uge_8131;
  reg p22_uge_8211;
  reg p22_uge_8291;
  reg [31:0] p22_concat_8370;
  reg p22_uge_8371;
  reg p22_bit_slice_6599;
  reg p22_bit_slice_6600;
  reg p22_bit_slice_6601;
  reg p22_bit_slice_6602;
  reg p22_bit_slice_6603;
  reg p22_bit_slice_6604;
  reg p22_bit_slice_6605;
  reg p22_bit_slice_6606;
  reg p22_bit_slice_6607;
  reg p22_negated;
  reg [31:0] p23_b;
  reg p23_uge_6683;
  reg [32:0] p23_bivisor__1;
  reg p23_uge_6691;
  reg p23_uge_6771;
  reg p23_uge_6851;
  reg p23_uge_6931;
  reg p23_uge_7011;
  reg p23_uge_7091;
  reg p23_uge_7171;
  reg p23_uge_7251;
  reg p23_uge_7331;
  reg p23_uge_7411;
  reg p23_uge_7491;
  reg p23_uge_7571;
  reg p23_uge_7651;
  reg p23_uge_7731;
  reg p23_uge_7811;
  reg p23_uge_7891;
  reg p23_uge_7971;
  reg p23_uge_8051;
  reg p23_uge_8131;
  reg p23_uge_8211;
  reg p23_uge_8291;
  reg p23_uge_8371;
  reg [31:0] p23_concat_8450;
  reg p23_uge_8451;
  reg p23_bit_slice_6600;
  reg p23_bit_slice_6601;
  reg p23_bit_slice_6602;
  reg p23_bit_slice_6603;
  reg p23_bit_slice_6604;
  reg p23_bit_slice_6605;
  reg p23_bit_slice_6606;
  reg p23_bit_slice_6607;
  reg p23_negated;
  reg [31:0] p24_b;
  reg p24_uge_6683;
  reg [32:0] p24_bivisor__1;
  reg p24_uge_6691;
  reg p24_uge_6771;
  reg p24_uge_6851;
  reg p24_uge_6931;
  reg p24_uge_7011;
  reg p24_uge_7091;
  reg p24_uge_7171;
  reg p24_uge_7251;
  reg p24_uge_7331;
  reg p24_uge_7411;
  reg p24_uge_7491;
  reg p24_uge_7571;
  reg p24_uge_7651;
  reg p24_uge_7731;
  reg p24_uge_7811;
  reg p24_uge_7891;
  reg p24_uge_7971;
  reg p24_uge_8051;
  reg p24_uge_8131;
  reg p24_uge_8211;
  reg p24_uge_8291;
  reg p24_uge_8371;
  reg p24_uge_8451;
  reg [31:0] p24_concat_8530;
  reg p24_uge_8531;
  reg p24_bit_slice_6601;
  reg p24_bit_slice_6602;
  reg p24_bit_slice_6603;
  reg p24_bit_slice_6604;
  reg p24_bit_slice_6605;
  reg p24_bit_slice_6606;
  reg p24_bit_slice_6607;
  reg p24_negated;
  reg [31:0] p25_b;
  reg p25_uge_6683;
  reg [32:0] p25_bivisor__1;
  reg p25_uge_6691;
  reg p25_uge_6771;
  reg p25_uge_6851;
  reg p25_uge_6931;
  reg p25_uge_7011;
  reg p25_uge_7091;
  reg p25_uge_7171;
  reg p25_uge_7251;
  reg p25_uge_7331;
  reg p25_uge_7411;
  reg p25_uge_7491;
  reg p25_uge_7571;
  reg p25_uge_7651;
  reg p25_uge_7731;
  reg p25_uge_7811;
  reg p25_uge_7891;
  reg p25_uge_7971;
  reg p25_uge_8051;
  reg p25_uge_8131;
  reg p25_uge_8211;
  reg p25_uge_8291;
  reg p25_uge_8371;
  reg p25_uge_8451;
  reg p25_uge_8531;
  reg [31:0] p25_concat_8610;
  reg p25_uge_8611;
  reg p25_bit_slice_6602;
  reg p25_bit_slice_6603;
  reg p25_bit_slice_6604;
  reg p25_bit_slice_6605;
  reg p25_bit_slice_6606;
  reg p25_bit_slice_6607;
  reg p25_negated;
  reg [31:0] p26_b;
  reg p26_uge_6683;
  reg [32:0] p26_bivisor__1;
  reg p26_uge_6691;
  reg p26_uge_6771;
  reg p26_uge_6851;
  reg p26_uge_6931;
  reg p26_uge_7011;
  reg p26_uge_7091;
  reg p26_uge_7171;
  reg p26_uge_7251;
  reg p26_uge_7331;
  reg p26_uge_7411;
  reg p26_uge_7491;
  reg p26_uge_7571;
  reg p26_uge_7651;
  reg p26_uge_7731;
  reg p26_uge_7811;
  reg p26_uge_7891;
  reg p26_uge_7971;
  reg p26_uge_8051;
  reg p26_uge_8131;
  reg p26_uge_8211;
  reg p26_uge_8291;
  reg p26_uge_8371;
  reg p26_uge_8451;
  reg p26_uge_8531;
  reg p26_uge_8611;
  reg [31:0] p26_concat_8690;
  reg p26_uge_8691;
  reg p26_bit_slice_6603;
  reg p26_bit_slice_6604;
  reg p26_bit_slice_6605;
  reg p26_bit_slice_6606;
  reg p26_bit_slice_6607;
  reg p26_negated;
  reg [31:0] p27_b;
  reg p27_uge_6683;
  reg [32:0] p27_bivisor__1;
  reg p27_uge_6691;
  reg p27_uge_6771;
  reg p27_uge_6851;
  reg p27_uge_6931;
  reg p27_uge_7011;
  reg p27_uge_7091;
  reg p27_uge_7171;
  reg p27_uge_7251;
  reg p27_uge_7331;
  reg p27_uge_7411;
  reg p27_uge_7491;
  reg p27_uge_7571;
  reg p27_uge_7651;
  reg p27_uge_7731;
  reg p27_uge_7811;
  reg p27_uge_7891;
  reg p27_uge_7971;
  reg p27_uge_8051;
  reg p27_uge_8131;
  reg p27_uge_8211;
  reg p27_uge_8291;
  reg p27_uge_8371;
  reg p27_uge_8451;
  reg p27_uge_8531;
  reg p27_uge_8611;
  reg p27_uge_8691;
  reg [31:0] p27_concat_8770;
  reg p27_uge_8771;
  reg p27_bit_slice_6604;
  reg p27_bit_slice_6605;
  reg p27_bit_slice_6606;
  reg p27_bit_slice_6607;
  reg p27_negated;
  reg [31:0] p28_b;
  reg p28_uge_6683;
  reg [32:0] p28_bivisor__1;
  reg p28_uge_6691;
  reg p28_uge_6771;
  reg p28_uge_6851;
  reg p28_uge_6931;
  reg p28_uge_7011;
  reg p28_uge_7091;
  reg p28_uge_7171;
  reg p28_uge_7251;
  reg p28_uge_7331;
  reg p28_uge_7411;
  reg p28_uge_7491;
  reg p28_uge_7571;
  reg p28_uge_7651;
  reg p28_uge_7731;
  reg p28_uge_7811;
  reg p28_uge_7891;
  reg p28_uge_7971;
  reg p28_uge_8051;
  reg p28_uge_8131;
  reg p28_uge_8211;
  reg p28_uge_8291;
  reg p28_uge_8371;
  reg p28_uge_8451;
  reg p28_uge_8531;
  reg p28_uge_8611;
  reg p28_uge_8691;
  reg p28_uge_8771;
  reg [31:0] p28_concat_8850;
  reg p28_uge_8851;
  reg p28_bit_slice_6605;
  reg p28_bit_slice_6606;
  reg p28_bit_slice_6607;
  reg p28_negated;
  reg [31:0] p29_b;
  reg p29_uge_6683;
  reg [32:0] p29_bivisor__1;
  reg p29_uge_6691;
  reg p29_uge_6771;
  reg p29_uge_6851;
  reg p29_uge_6931;
  reg p29_uge_7011;
  reg p29_uge_7091;
  reg p29_uge_7171;
  reg p29_uge_7251;
  reg p29_uge_7331;
  reg p29_uge_7411;
  reg p29_uge_7491;
  reg p29_uge_7571;
  reg p29_uge_7651;
  reg p29_uge_7731;
  reg p29_uge_7811;
  reg p29_uge_7891;
  reg p29_uge_7971;
  reg p29_uge_8051;
  reg p29_uge_8131;
  reg p29_uge_8211;
  reg p29_uge_8291;
  reg p29_uge_8371;
  reg p29_uge_8451;
  reg p29_uge_8531;
  reg p29_uge_8611;
  reg p29_uge_8691;
  reg p29_uge_8771;
  reg p29_uge_8851;
  reg [31:0] p29_concat_8930;
  reg p29_uge_8931;
  reg p29_bit_slice_6606;
  reg p29_bit_slice_6607;
  reg p29_negated;
  reg [31:0] p30_b;
  reg p30_uge_6683;
  reg [32:0] p30_bivisor__1;
  reg p30_uge_6691;
  reg p30_uge_6771;
  reg p30_uge_6851;
  reg p30_uge_6931;
  reg p30_uge_7011;
  reg p30_uge_7091;
  reg p30_uge_7171;
  reg p30_uge_7251;
  reg p30_uge_7331;
  reg p30_uge_7411;
  reg p30_uge_7491;
  reg p30_uge_7571;
  reg p30_uge_7651;
  reg p30_uge_7731;
  reg p30_uge_7811;
  reg p30_uge_7891;
  reg p30_uge_7971;
  reg p30_uge_8051;
  reg p30_uge_8131;
  reg p30_uge_8211;
  reg p30_uge_8291;
  reg p30_uge_8371;
  reg p30_uge_8451;
  reg p30_uge_8531;
  reg p30_uge_8611;
  reg p30_uge_8691;
  reg p30_uge_8771;
  reg p30_uge_8851;
  reg p30_uge_8931;
  reg [31:0] p30_concat_9010;
  reg p30_uge_9011;
  reg p30_bit_slice_6607;
  reg p30_negated;
  reg p31_uge_6683;
  reg p31_uge_6691;
  reg p31_uge_6771;
  reg p31_uge_6851;
  reg p31_uge_6931;
  reg p31_uge_7011;
  reg p31_uge_7091;
  reg p31_uge_7171;
  reg p31_uge_7251;
  reg p31_uge_7331;
  reg p31_uge_7411;
  reg p31_uge_7491;
  reg p31_uge_7571;
  reg p31_uge_7651;
  reg p31_uge_7731;
  reg p31_uge_7811;
  reg p31_uge_7891;
  reg p31_uge_7971;
  reg p31_uge_8051;
  reg p31_uge_8131;
  reg p31_uge_8211;
  reg p31_uge_8291;
  reg p31_uge_8371;
  reg p31_uge_8451;
  reg p31_uge_8531;
  reg p31_uge_8611;
  reg p31_uge_8691;
  reg p31_uge_8771;
  reg p31_uge_8851;
  reg p31_uge_8931;
  reg p31_uge_9011;
  reg p31_q__32_squeezed_portion_0_width_1;
  reg p31_negated;
  reg p0_valid;
  reg p1_valid;
  reg p2_valid;
  reg p3_valid;
  reg p4_valid;
  reg p5_valid;
  reg p6_valid;
  reg p7_valid;
  reg p8_valid;
  reg p9_valid;
  reg p10_valid;
  reg p11_valid;
  reg p12_valid;
  reg p13_valid;
  reg p14_valid;
  reg p15_valid;
  reg p16_valid;
  reg p17_valid;
  reg p18_valid;
  reg p19_valid;
  reg p20_valid;
  reg p21_valid;
  reg p22_valid;
  reg p23_valid;
  reg p24_valid;
  reg p25_valid;
  reg p26_valid;
  reg p27_valid;
  reg p28_valid;
  reg p29_valid;
  reg p30_valid;
  reg p31_valid;
  reg p32_valid;
  reg p33_valid;
  reg p34_valid;
  reg [31:0] __xls_float_ips__result_reg;
  reg __xls_float_ips__result_valid_reg;
  wire xls_float_ips__result_valid_inv;
  wire xls_float_ips__result_valid_load_en;
  wire xls_float_ips__result_load_en;
  wire p32_stage_done;
  wire p32_not_valid;
  wire p31_enable;
  wire p31_data_enable;
  wire p31_not_valid;
  wire p30_enable;
  wire p30_data_enable;
  wire p30_not_valid;
  wire p29_enable;
  wire p29_data_enable;
  wire p29_not_valid;
  wire p28_enable;
  wire p28_data_enable;
  wire p28_not_valid;
  wire p27_enable;
  wire p27_data_enable;
  wire p27_not_valid;
  wire p26_enable;
  wire p26_data_enable;
  wire p26_not_valid;
  wire p25_enable;
  wire p25_data_enable;
  wire p25_not_valid;
  wire p24_enable;
  wire p24_data_enable;
  wire p24_not_valid;
  wire p23_enable;
  wire p23_data_enable;
  wire p23_not_valid;
  wire p22_enable;
  wire p22_data_enable;
  wire p22_not_valid;
  wire p21_enable;
  wire p21_data_enable;
  wire p21_not_valid;
  wire p20_enable;
  wire p20_data_enable;
  wire p20_not_valid;
  wire p19_enable;
  wire p19_data_enable;
  wire p19_not_valid;
  wire p18_enable;
  wire p18_data_enable;
  wire p18_not_valid;
  wire p17_enable;
  wire p17_data_enable;
  wire p17_not_valid;
  wire p16_enable;
  wire p16_data_enable;
  wire p16_not_valid;
  wire p15_enable;
  wire p15_data_enable;
  wire p15_not_valid;
  wire p14_enable;
  wire p14_data_enable;
  wire p14_not_valid;
  wire p13_enable;
  wire p13_data_enable;
  wire p13_not_valid;
  wire p12_enable;
  wire p12_data_enable;
  wire p12_not_valid;
  wire p11_enable;
  wire p11_data_enable;
  wire p11_not_valid;
  wire p10_enable;
  wire p10_data_enable;
  wire p10_not_valid;
  wire p9_enable;
  wire p9_data_enable;
  wire p9_not_valid;
  wire p8_enable;
  wire p8_data_enable;
  wire p8_not_valid;
  wire p7_enable;
  wire p7_data_enable;
  wire p7_not_valid;
  wire p6_enable;
  wire p6_data_enable;
  wire p6_not_valid;
  wire p5_enable;
  wire p5_data_enable;
  wire p5_not_valid;
  wire p4_enable;
  wire p4_data_enable;
  wire p4_not_valid;
  wire p3_enable;
  wire p3_data_enable;
  wire p3_not_valid;
  wire p2_enable;
  wire p2_data_enable;
  wire p2_not_valid;
  wire [31:0] sub_9086;
  wire [31:0] sub_9006;
  wire [31:0] sub_8926;
  wire [31:0] sub_8846;
  wire [31:0] sub_8766;
  wire [31:0] sub_8686;
  wire [31:0] sub_8606;
  wire [31:0] sub_8526;
  wire [31:0] sub_8446;
  wire [31:0] sub_8366;
  wire [31:0] sub_8286;
  wire [31:0] sub_8206;
  wire [31:0] sub_8126;
  wire [31:0] sub_8046;
  wire [31:0] sub_7966;
  wire [31:0] sub_7886;
  wire [31:0] sub_7806;
  wire [31:0] sub_7726;
  wire [31:0] sub_7646;
  wire [31:0] sub_7566;
  wire [31:0] sub_7486;
  wire [31:0] sub_7406;
  wire [31:0] sub_7326;
  wire [31:0] sub_7246;
  wire [31:0] sub_7166;
  wire [31:0] sub_7086;
  wire [31:0] sub_7006;
  wire [31:0] sub_6926;
  wire [31:0] sub_6846;
  wire [31:0] sub_6766;
  wire uge_6683;
  wire [31:0] sub_6684;
  wire p1_enable;
  wire [31:0] r__62;
  wire [31:0] r__60;
  wire [31:0] r__58;
  wire [31:0] r__56;
  wire [31:0] r__54;
  wire [31:0] r__52;
  wire [31:0] r__50;
  wire [31:0] r__48;
  wire [31:0] r__46;
  wire [31:0] r__44;
  wire [31:0] r__42;
  wire [31:0] r__40;
  wire [31:0] r__38;
  wire [31:0] r__36;
  wire [31:0] r__34;
  wire [31:0] r__32;
  wire [31:0] r__30;
  wire [31:0] r__28;
  wire [31:0] r__26;
  wire [31:0] r__24;
  wire [31:0] r__22;
  wire [31:0] r__20;
  wire [31:0] r__18;
  wire [31:0] r__16;
  wire [31:0] r__14;
  wire [31:0] r__12;
  wire [31:0] r__10;
  wire [31:0] r__8;
  wire [31:0] r__6;
  wire [31:0] r__4;
  wire [31:0] r__2;
  wire p1_data_enable;
  wire p1_not_valid;
  wire [31:0] q__32;
  wire [32:0] r__63;
  wire [32:0] r__61;
  wire [32:0] r__59;
  wire [32:0] r__57;
  wire [32:0] r__55;
  wire [32:0] r__53;
  wire [32:0] r__51;
  wire [32:0] r__49;
  wire [32:0] r__47;
  wire [32:0] r__45;
  wire [32:0] r__43;
  wire [32:0] r__41;
  wire [32:0] r__39;
  wire [32:0] r__37;
  wire [32:0] r__35;
  wire [32:0] r__33;
  wire [32:0] r__31;
  wire [32:0] r__29;
  wire [32:0] r__27;
  wire [32:0] r__25;
  wire [32:0] r__23;
  wire [32:0] r__21;
  wire [32:0] r__19;
  wire [32:0] r__17;
  wire [32:0] r__15;
  wire [32:0] r__13;
  wire [32:0] r__11;
  wire [32:0] r__9;
  wire [32:0] r__7;
  wire [32:0] r__5;
  wire [32:0] r__3;
  wire [32:0] bivisor__1;
  wire sign_a;
  wire p0_enable;
  wire p0_all_active_inputs_valid;
  wire sign_b;
  wire p34_enable;
  wire p33_enable;
  wire p32_enable;
  wire q__32_squeezed_portion_0_width_1;
  wire [31:0] concat_9010;
  wire uge_9011;
  wire [31:0] concat_8930;
  wire uge_8931;
  wire [31:0] concat_8850;
  wire uge_8851;
  wire [31:0] concat_8770;
  wire uge_8771;
  wire [31:0] concat_8690;
  wire uge_8691;
  wire [31:0] concat_8610;
  wire uge_8611;
  wire [31:0] concat_8530;
  wire uge_8531;
  wire [31:0] concat_8450;
  wire uge_8451;
  wire [31:0] concat_8370;
  wire uge_8371;
  wire [31:0] concat_8290;
  wire uge_8291;
  wire [31:0] concat_8210;
  wire uge_8211;
  wire [31:0] concat_8130;
  wire uge_8131;
  wire [31:0] concat_8050;
  wire uge_8051;
  wire [31:0] concat_7970;
  wire uge_7971;
  wire [31:0] concat_7890;
  wire uge_7891;
  wire [31:0] concat_7810;
  wire uge_7811;
  wire [31:0] concat_7730;
  wire uge_7731;
  wire [31:0] concat_7650;
  wire uge_7651;
  wire [31:0] concat_7570;
  wire uge_7571;
  wire [31:0] concat_7490;
  wire uge_7491;
  wire [31:0] concat_7410;
  wire uge_7411;
  wire [31:0] concat_7330;
  wire uge_7331;
  wire [31:0] concat_7250;
  wire uge_7251;
  wire [31:0] concat_7170;
  wire uge_7171;
  wire [31:0] concat_7090;
  wire uge_7091;
  wire [31:0] concat_7010;
  wire uge_7011;
  wire [31:0] concat_6930;
  wire uge_6931;
  wire [31:0] concat_6850;
  wire uge_6851;
  wire [31:0] concat_6770;
  wire uge_6771;
  wire [31:0] concat_6690;
  wire uge_6691;
  wire [31:0] concat_6575;
  wire p0_data_enable;
  wire bit_slice_6577;
  wire bit_slice_6578;
  wire bit_slice_6579;
  wire bit_slice_6580;
  wire bit_slice_6581;
  wire bit_slice_6582;
  wire bit_slice_6583;
  wire bit_slice_6584;
  wire bit_slice_6585;
  wire bit_slice_6586;
  wire bit_slice_6587;
  wire bit_slice_6588;
  wire bit_slice_6589;
  wire bit_slice_6590;
  wire bit_slice_6591;
  wire bit_slice_6592;
  wire bit_slice_6593;
  wire bit_slice_6594;
  wire bit_slice_6595;
  wire bit_slice_6596;
  wire bit_slice_6597;
  wire bit_slice_6598;
  wire bit_slice_6599;
  wire bit_slice_6600;
  wire bit_slice_6601;
  wire bit_slice_6602;
  wire bit_slice_6603;
  wire bit_slice_6604;
  wire bit_slice_6605;
  wire bit_slice_6606;
  wire bit_slice_6607;
  wire negated;
  wire [31:0] __xls_float_ips__result_buf;
  assign xls_float_ips__result_valid_inv = ~__xls_float_ips__result_valid_reg;
  assign xls_float_ips__result_valid_load_en = xls_float_ips__result_rdy | xls_float_ips__result_valid_inv;
  assign xls_float_ips__result_load_en = p31_valid & xls_float_ips__result_valid_load_en;
  assign p32_stage_done = p31_valid & xls_float_ips__result_load_en;
  assign p32_not_valid = ~p31_valid;
  assign p31_enable = p32_stage_done | p32_not_valid;
  assign p31_data_enable = p31_enable & p30_valid;
  assign p31_not_valid = ~p30_valid;
  assign p30_enable = p31_data_enable | p31_not_valid;
  assign p30_data_enable = p30_enable & p29_valid;
  assign p30_not_valid = ~p29_valid;
  assign p29_enable = p30_data_enable | p30_not_valid;
  assign p29_data_enable = p29_enable & p28_valid;
  assign p29_not_valid = ~p28_valid;
  assign p28_enable = p29_data_enable | p29_not_valid;
  assign p28_data_enable = p28_enable & p27_valid;
  assign p28_not_valid = ~p27_valid;
  assign p27_enable = p28_data_enable | p28_not_valid;
  assign p27_data_enable = p27_enable & p26_valid;
  assign p27_not_valid = ~p26_valid;
  assign p26_enable = p27_data_enable | p27_not_valid;
  assign p26_data_enable = p26_enable & p25_valid;
  assign p26_not_valid = ~p25_valid;
  assign p25_enable = p26_data_enable | p26_not_valid;
  assign p25_data_enable = p25_enable & p24_valid;
  assign p25_not_valid = ~p24_valid;
  assign p24_enable = p25_data_enable | p25_not_valid;
  assign p24_data_enable = p24_enable & p23_valid;
  assign p24_not_valid = ~p23_valid;
  assign p23_enable = p24_data_enable | p24_not_valid;
  assign p23_data_enable = p23_enable & p22_valid;
  assign p23_not_valid = ~p22_valid;
  assign p22_enable = p23_data_enable | p23_not_valid;
  assign p22_data_enable = p22_enable & p21_valid;
  assign p22_not_valid = ~p21_valid;
  assign p21_enable = p22_data_enable | p22_not_valid;
  assign p21_data_enable = p21_enable & p20_valid;
  assign p21_not_valid = ~p20_valid;
  assign p20_enable = p21_data_enable | p21_not_valid;
  assign p20_data_enable = p20_enable & p19_valid;
  assign p20_not_valid = ~p19_valid;
  assign p19_enable = p20_data_enable | p20_not_valid;
  assign p19_data_enable = p19_enable & p18_valid;
  assign p19_not_valid = ~p18_valid;
  assign p18_enable = p19_data_enable | p19_not_valid;
  assign p18_data_enable = p18_enable & p17_valid;
  assign p18_not_valid = ~p17_valid;
  assign p17_enable = p18_data_enable | p18_not_valid;
  assign p17_data_enable = p17_enable & p16_valid;
  assign p17_not_valid = ~p16_valid;
  assign p16_enable = p17_data_enable | p17_not_valid;
  assign p16_data_enable = p16_enable & p15_valid;
  assign p16_not_valid = ~p15_valid;
  assign p15_enable = p16_data_enable | p16_not_valid;
  assign p15_data_enable = p15_enable & p14_valid;
  assign p15_not_valid = ~p14_valid;
  assign p14_enable = p15_data_enable | p15_not_valid;
  assign p14_data_enable = p14_enable & p13_valid;
  assign p14_not_valid = ~p13_valid;
  assign p13_enable = p14_data_enable | p14_not_valid;
  assign p13_data_enable = p13_enable & p12_valid;
  assign p13_not_valid = ~p12_valid;
  assign p12_enable = p13_data_enable | p13_not_valid;
  assign p12_data_enable = p12_enable & p11_valid;
  assign p12_not_valid = ~p11_valid;
  assign p11_enable = p12_data_enable | p12_not_valid;
  assign p11_data_enable = p11_enable & p10_valid;
  assign p11_not_valid = ~p10_valid;
  assign p10_enable = p11_data_enable | p11_not_valid;
  assign p10_data_enable = p10_enable & p9_valid;
  assign p10_not_valid = ~p9_valid;
  assign p9_enable = p10_data_enable | p10_not_valid;
  assign p9_data_enable = p9_enable & p8_valid;
  assign p9_not_valid = ~p8_valid;
  assign p8_enable = p9_data_enable | p9_not_valid;
  assign p8_data_enable = p8_enable & p7_valid;
  assign p8_not_valid = ~p7_valid;
  assign p7_enable = p8_data_enable | p8_not_valid;
  assign p7_data_enable = p7_enable & p6_valid;
  assign p7_not_valid = ~p6_valid;
  assign p6_enable = p7_data_enable | p7_not_valid;
  assign p6_data_enable = p6_enable & p5_valid;
  assign p6_not_valid = ~p5_valid;
  assign p5_enable = p6_data_enable | p6_not_valid;
  assign p5_data_enable = p5_enable & p4_valid;
  assign p5_not_valid = ~p4_valid;
  assign p4_enable = p5_data_enable | p5_not_valid;
  assign p4_data_enable = p4_enable & p3_valid;
  assign p4_not_valid = ~p3_valid;
  assign p3_enable = p4_data_enable | p4_not_valid;
  assign p3_data_enable = p3_enable & p2_valid;
  assign p3_not_valid = ~p2_valid;
  assign p2_enable = p3_data_enable | p3_not_valid;
  assign p2_data_enable = p2_enable & p1_valid;
  assign p2_not_valid = ~p1_valid;
  assign sub_9086 = p30_concat_9010 - p30_b;
  assign sub_9006 = p29_concat_8930 - p29_b;
  assign sub_8926 = p28_concat_8850 - p28_b;
  assign sub_8846 = p27_concat_8770 - p27_b;
  assign sub_8766 = p26_concat_8690 - p26_b;
  assign sub_8686 = p25_concat_8610 - p25_b;
  assign sub_8606 = p24_concat_8530 - p24_b;
  assign sub_8526 = p23_concat_8450 - p23_b;
  assign sub_8446 = p22_concat_8370 - p22_b;
  assign sub_8366 = p21_concat_8290 - p21_b;
  assign sub_8286 = p20_concat_8210 - p20_b;
  assign sub_8206 = p19_concat_8130 - p19_b;
  assign sub_8126 = p18_concat_8050 - p18_b;
  assign sub_8046 = p17_concat_7970 - p17_b;
  assign sub_7966 = p16_concat_7890 - p16_b;
  assign sub_7886 = p15_concat_7810 - p15_b;
  assign sub_7806 = p14_concat_7730 - p14_b;
  assign sub_7726 = p13_concat_7650 - p13_b;
  assign sub_7646 = p12_concat_7570 - p12_b;
  assign sub_7566 = p11_concat_7490 - p11_b;
  assign sub_7486 = p10_concat_7410 - p10_b;
  assign sub_7406 = p9_concat_7330 - p9_b;
  assign sub_7326 = p8_concat_7250 - p8_b;
  assign sub_7246 = p7_concat_7170 - p7_b;
  assign sub_7166 = p6_concat_7090 - p6_b;
  assign sub_7086 = p5_concat_7010 - p5_b;
  assign sub_7006 = p4_concat_6930 - p4_b;
  assign sub_6926 = p3_concat_6850 - p3_b;
  assign sub_6846 = p2_concat_6770 - p2_b;
  assign sub_6766 = p1_concat_6690 - p1_b;
  assign uge_6683 = p0_concat_6575 >= p0_b;
  assign sub_6684 = p0_concat_6575 - p0_b;
  assign p1_enable = p2_data_enable | p2_not_valid;
  assign r__62 = p30_uge_9011 ? sub_9086 : p30_concat_9010;
  assign r__60 = p29_uge_8931 ? sub_9006 : p29_concat_8930;
  assign r__58 = p28_uge_8851 ? sub_8926 : p28_concat_8850;
  assign r__56 = p27_uge_8771 ? sub_8846 : p27_concat_8770;
  assign r__54 = p26_uge_8691 ? sub_8766 : p26_concat_8690;
  assign r__52 = p25_uge_8611 ? sub_8686 : p25_concat_8610;
  assign r__50 = p24_uge_8531 ? sub_8606 : p24_concat_8530;
  assign r__48 = p23_uge_8451 ? sub_8526 : p23_concat_8450;
  assign r__46 = p22_uge_8371 ? sub_8446 : p22_concat_8370;
  assign r__44 = p21_uge_8291 ? sub_8366 : p21_concat_8290;
  assign r__42 = p20_uge_8211 ? sub_8286 : p20_concat_8210;
  assign r__40 = p19_uge_8131 ? sub_8206 : p19_concat_8130;
  assign r__38 = p18_uge_8051 ? sub_8126 : p18_concat_8050;
  assign r__36 = p17_uge_7971 ? sub_8046 : p17_concat_7970;
  assign r__34 = p16_uge_7891 ? sub_7966 : p16_concat_7890;
  assign r__32 = p15_uge_7811 ? sub_7886 : p15_concat_7810;
  assign r__30 = p14_uge_7731 ? sub_7806 : p14_concat_7730;
  assign r__28 = p13_uge_7651 ? sub_7726 : p13_concat_7650;
  assign r__26 = p12_uge_7571 ? sub_7646 : p12_concat_7570;
  assign r__24 = p11_uge_7491 ? sub_7566 : p11_concat_7490;
  assign r__22 = p10_uge_7411 ? sub_7486 : p10_concat_7410;
  assign r__20 = p9_uge_7331 ? sub_7406 : p9_concat_7330;
  assign r__18 = p8_uge_7251 ? sub_7326 : p8_concat_7250;
  assign r__16 = p7_uge_7171 ? sub_7246 : p7_concat_7170;
  assign r__14 = p6_uge_7091 ? sub_7166 : p6_concat_7090;
  assign r__12 = p5_uge_7011 ? sub_7086 : p5_concat_7010;
  assign r__10 = p4_uge_6931 ? sub_7006 : p4_concat_6930;
  assign r__8 = p3_uge_6851 ? sub_6926 : p3_concat_6850;
  assign r__6 = p2_uge_6771 ? sub_6846 : p2_concat_6770;
  assign r__4 = p1_uge_6691 ? sub_6766 : p1_concat_6690;
  assign r__2 = uge_6683 ? sub_6684 : p0_concat_6575;
  assign p1_data_enable = p1_enable & p0_valid;
  assign p1_not_valid = ~p0_valid;
  assign q__32 = {p31_uge_6683, p31_uge_6691, p31_uge_6771, p31_uge_6851, p31_uge_6931, p31_uge_7011, p31_uge_7091, p31_uge_7171, p31_uge_7251, p31_uge_7331, p31_uge_7411, p31_uge_7491, p31_uge_7571, p31_uge_7651, p31_uge_7731, p31_uge_7811, p31_uge_7891, p31_uge_7971, p31_uge_8051, p31_uge_8131, p31_uge_8211, p31_uge_8291, p31_uge_8371, p31_uge_8451, p31_uge_8531, p31_uge_8611, p31_uge_8691, p31_uge_8771, p31_uge_8851, p31_uge_8931, p31_uge_9011, p31_q__32_squeezed_portion_0_width_1};
  assign r__63 = {r__62, p30_bit_slice_6607};
  assign r__61 = {r__60, p29_bit_slice_6606};
  assign r__59 = {r__58, p28_bit_slice_6605};
  assign r__57 = {r__56, p27_bit_slice_6604};
  assign r__55 = {r__54, p26_bit_slice_6603};
  assign r__53 = {r__52, p25_bit_slice_6602};
  assign r__51 = {r__50, p24_bit_slice_6601};
  assign r__49 = {r__48, p23_bit_slice_6600};
  assign r__47 = {r__46, p22_bit_slice_6599};
  assign r__45 = {r__44, p21_bit_slice_6598};
  assign r__43 = {r__42, p20_bit_slice_6597};
  assign r__41 = {r__40, p19_bit_slice_6596};
  assign r__39 = {r__38, p18_bit_slice_6595};
  assign r__37 = {r__36, p17_bit_slice_6594};
  assign r__35 = {r__34, p16_bit_slice_6593};
  assign r__33 = {r__32, p15_bit_slice_6592};
  assign r__31 = {r__30, p14_bit_slice_6591};
  assign r__29 = {r__28, p13_bit_slice_6590};
  assign r__27 = {r__26, p12_bit_slice_6589};
  assign r__25 = {r__24, p11_bit_slice_6588};
  assign r__23 = {r__22, p10_bit_slice_6587};
  assign r__21 = {r__20, p9_bit_slice_6586};
  assign r__19 = {r__18, p8_bit_slice_6585};
  assign r__17 = {r__16, p7_bit_slice_6584};
  assign r__15 = {r__14, p6_bit_slice_6583};
  assign r__13 = {r__12, p5_bit_slice_6582};
  assign r__11 = {r__10, p4_bit_slice_6581};
  assign r__9 = {r__8, p3_bit_slice_6580};
  assign r__7 = {r__6, p2_bit_slice_6579};
  assign r__5 = {r__4, p1_bit_slice_6578};
  assign r__3 = {r__2, p0_bit_slice_6577};
  assign bivisor__1 = {1'h0, p0_b};
  assign sign_a = xls_float_ips__lhs[31];
  assign p0_enable = p1_data_enable | p1_not_valid;
  assign p0_all_active_inputs_valid = xls_float_ips__lhs_vld & xls_float_ips__rhs_vld;
  assign sign_b = xls_float_ips__rhs[31];
  assign p34_enable = 1'h1;
  assign p33_enable = 1'h1;
  assign p32_enable = 1'h1;
  assign q__32_squeezed_portion_0_width_1 = r__63 >= p30_bivisor__1;
  assign concat_9010 = {r__60[30:0], p29_bit_slice_6606};
  assign uge_9011 = r__61 >= p29_bivisor__1;
  assign concat_8930 = {r__58[30:0], p28_bit_slice_6605};
  assign uge_8931 = r__59 >= p28_bivisor__1;
  assign concat_8850 = {r__56[30:0], p27_bit_slice_6604};
  assign uge_8851 = r__57 >= p27_bivisor__1;
  assign concat_8770 = {r__54[30:0], p26_bit_slice_6603};
  assign uge_8771 = r__55 >= p26_bivisor__1;
  assign concat_8690 = {r__52[30:0], p25_bit_slice_6602};
  assign uge_8691 = r__53 >= p25_bivisor__1;
  assign concat_8610 = {r__50[30:0], p24_bit_slice_6601};
  assign uge_8611 = r__51 >= p24_bivisor__1;
  assign concat_8530 = {r__48[30:0], p23_bit_slice_6600};
  assign uge_8531 = r__49 >= p23_bivisor__1;
  assign concat_8450 = {r__46[30:0], p22_bit_slice_6599};
  assign uge_8451 = r__47 >= p22_bivisor__1;
  assign concat_8370 = {r__44[30:0], p21_bit_slice_6598};
  assign uge_8371 = r__45 >= p21_bivisor__1;
  assign concat_8290 = {r__42[30:0], p20_bit_slice_6597};
  assign uge_8291 = r__43 >= p20_bivisor__1;
  assign concat_8210 = {r__40[30:0], p19_bit_slice_6596};
  assign uge_8211 = r__41 >= p19_bivisor__1;
  assign concat_8130 = {r__38[30:0], p18_bit_slice_6595};
  assign uge_8131 = r__39 >= p18_bivisor__1;
  assign concat_8050 = {r__36[30:0], p17_bit_slice_6594};
  assign uge_8051 = r__37 >= p17_bivisor__1;
  assign concat_7970 = {r__34[30:0], p16_bit_slice_6593};
  assign uge_7971 = r__35 >= p16_bivisor__1;
  assign concat_7890 = {r__32[30:0], p15_bit_slice_6592};
  assign uge_7891 = r__33 >= p15_bivisor__1;
  assign concat_7810 = {r__30[30:0], p14_bit_slice_6591};
  assign uge_7811 = r__31 >= p14_bivisor__1;
  assign concat_7730 = {r__28[30:0], p13_bit_slice_6590};
  assign uge_7731 = r__29 >= p13_bivisor__1;
  assign concat_7650 = {r__26[30:0], p12_bit_slice_6589};
  assign uge_7651 = r__27 >= p12_bivisor__1;
  assign concat_7570 = {r__24[30:0], p11_bit_slice_6588};
  assign uge_7571 = r__25 >= p11_bivisor__1;
  assign concat_7490 = {r__22[30:0], p10_bit_slice_6587};
  assign uge_7491 = r__23 >= p10_bivisor__1;
  assign concat_7410 = {r__20[30:0], p9_bit_slice_6586};
  assign uge_7411 = r__21 >= p9_bivisor__1;
  assign concat_7330 = {r__18[30:0], p8_bit_slice_6585};
  assign uge_7331 = r__19 >= p8_bivisor__1;
  assign concat_7250 = {r__16[30:0], p7_bit_slice_6584};
  assign uge_7251 = r__17 >= p7_bivisor__1;
  assign concat_7170 = {r__14[30:0], p6_bit_slice_6583};
  assign uge_7171 = r__15 >= p6_bivisor__1;
  assign concat_7090 = {r__12[30:0], p5_bit_slice_6582};
  assign uge_7091 = r__13 >= p5_bivisor__1;
  assign concat_7010 = {r__10[30:0], p4_bit_slice_6581};
  assign uge_7011 = r__11 >= p4_bivisor__1;
  assign concat_6930 = {r__8[30:0], p3_bit_slice_6580};
  assign uge_6931 = r__9 >= p3_bivisor__1;
  assign concat_6850 = {r__6[30:0], p2_bit_slice_6579};
  assign uge_6851 = r__7 >= p2_bivisor__1;
  assign concat_6770 = {r__4[30:0], p1_bit_slice_6578};
  assign uge_6771 = r__5 >= p1_bivisor__1;
  assign concat_6690 = {r__2[30:0], p0_bit_slice_6577};
  assign uge_6691 = r__3 >= bivisor__1;
  assign concat_6575 = {31'h0000_0000, sign_a};
  assign p0_data_enable = p0_enable & p0_all_active_inputs_valid;
  assign bit_slice_6577 = xls_float_ips__lhs[30];
  assign bit_slice_6578 = xls_float_ips__lhs[29];
  assign bit_slice_6579 = xls_float_ips__lhs[28];
  assign bit_slice_6580 = xls_float_ips__lhs[27];
  assign bit_slice_6581 = xls_float_ips__lhs[26];
  assign bit_slice_6582 = xls_float_ips__lhs[25];
  assign bit_slice_6583 = xls_float_ips__lhs[24];
  assign bit_slice_6584 = xls_float_ips__lhs[23];
  assign bit_slice_6585 = xls_float_ips__lhs[22];
  assign bit_slice_6586 = xls_float_ips__lhs[21];
  assign bit_slice_6587 = xls_float_ips__lhs[20];
  assign bit_slice_6588 = xls_float_ips__lhs[19];
  assign bit_slice_6589 = xls_float_ips__lhs[18];
  assign bit_slice_6590 = xls_float_ips__lhs[17];
  assign bit_slice_6591 = xls_float_ips__lhs[16];
  assign bit_slice_6592 = xls_float_ips__lhs[15];
  assign bit_slice_6593 = xls_float_ips__lhs[14];
  assign bit_slice_6594 = xls_float_ips__lhs[13];
  assign bit_slice_6595 = xls_float_ips__lhs[12];
  assign bit_slice_6596 = xls_float_ips__lhs[11];
  assign bit_slice_6597 = xls_float_ips__lhs[10];
  assign bit_slice_6598 = xls_float_ips__lhs[9];
  assign bit_slice_6599 = xls_float_ips__lhs[8];
  assign bit_slice_6600 = xls_float_ips__lhs[7];
  assign bit_slice_6601 = xls_float_ips__lhs[6];
  assign bit_slice_6602 = xls_float_ips__lhs[5];
  assign bit_slice_6603 = xls_float_ips__lhs[4];
  assign bit_slice_6604 = xls_float_ips__lhs[3];
  assign bit_slice_6605 = xls_float_ips__lhs[2];
  assign bit_slice_6606 = xls_float_ips__lhs[1];
  assign bit_slice_6607 = xls_float_ips__lhs[0];
  assign negated = sign_a ^ sign_b;
  assign __xls_float_ips__result_buf = p31_negated ? -q__32 : q__32;
  always @ (posedge clk) begin
    if (rst) begin
      p0_concat_6575 <= 32'h0000_0000;
      p0_b <= 32'h0000_0000;
      p0_bit_slice_6577 <= 1'h0;
      p0_bit_slice_6578 <= 1'h0;
      p0_bit_slice_6579 <= 1'h0;
      p0_bit_slice_6580 <= 1'h0;
      p0_bit_slice_6581 <= 1'h0;
      p0_bit_slice_6582 <= 1'h0;
      p0_bit_slice_6583 <= 1'h0;
      p0_bit_slice_6584 <= 1'h0;
      p0_bit_slice_6585 <= 1'h0;
      p0_bit_slice_6586 <= 1'h0;
      p0_bit_slice_6587 <= 1'h0;
      p0_bit_slice_6588 <= 1'h0;
      p0_bit_slice_6589 <= 1'h0;
      p0_bit_slice_6590 <= 1'h0;
      p0_bit_slice_6591 <= 1'h0;
      p0_bit_slice_6592 <= 1'h0;
      p0_bit_slice_6593 <= 1'h0;
      p0_bit_slice_6594 <= 1'h0;
      p0_bit_slice_6595 <= 1'h0;
      p0_bit_slice_6596 <= 1'h0;
      p0_bit_slice_6597 <= 1'h0;
      p0_bit_slice_6598 <= 1'h0;
      p0_bit_slice_6599 <= 1'h0;
      p0_bit_slice_6600 <= 1'h0;
      p0_bit_slice_6601 <= 1'h0;
      p0_bit_slice_6602 <= 1'h0;
      p0_bit_slice_6603 <= 1'h0;
      p0_bit_slice_6604 <= 1'h0;
      p0_bit_slice_6605 <= 1'h0;
      p0_bit_slice_6606 <= 1'h0;
      p0_bit_slice_6607 <= 1'h0;
      p0_negated <= 1'h0;
      p1_b <= 32'h0000_0000;
      p1_uge_6683 <= 1'h0;
      p1_bivisor__1 <= 33'h0_0000_0000;
      p1_concat_6690 <= 32'h0000_0000;
      p1_uge_6691 <= 1'h0;
      p1_bit_slice_6578 <= 1'h0;
      p1_bit_slice_6579 <= 1'h0;
      p1_bit_slice_6580 <= 1'h0;
      p1_bit_slice_6581 <= 1'h0;
      p1_bit_slice_6582 <= 1'h0;
      p1_bit_slice_6583 <= 1'h0;
      p1_bit_slice_6584 <= 1'h0;
      p1_bit_slice_6585 <= 1'h0;
      p1_bit_slice_6586 <= 1'h0;
      p1_bit_slice_6587 <= 1'h0;
      p1_bit_slice_6588 <= 1'h0;
      p1_bit_slice_6589 <= 1'h0;
      p1_bit_slice_6590 <= 1'h0;
      p1_bit_slice_6591 <= 1'h0;
      p1_bit_slice_6592 <= 1'h0;
      p1_bit_slice_6593 <= 1'h0;
      p1_bit_slice_6594 <= 1'h0;
      p1_bit_slice_6595 <= 1'h0;
      p1_bit_slice_6596 <= 1'h0;
      p1_bit_slice_6597 <= 1'h0;
      p1_bit_slice_6598 <= 1'h0;
      p1_bit_slice_6599 <= 1'h0;
      p1_bit_slice_6600 <= 1'h0;
      p1_bit_slice_6601 <= 1'h0;
      p1_bit_slice_6602 <= 1'h0;
      p1_bit_slice_6603 <= 1'h0;
      p1_bit_slice_6604 <= 1'h0;
      p1_bit_slice_6605 <= 1'h0;
      p1_bit_slice_6606 <= 1'h0;
      p1_bit_slice_6607 <= 1'h0;
      p1_negated <= 1'h0;
      p2_b <= 32'h0000_0000;
      p2_uge_6683 <= 1'h0;
      p2_bivisor__1 <= 33'h0_0000_0000;
      p2_uge_6691 <= 1'h0;
      p2_concat_6770 <= 32'h0000_0000;
      p2_uge_6771 <= 1'h0;
      p2_bit_slice_6579 <= 1'h0;
      p2_bit_slice_6580 <= 1'h0;
      p2_bit_slice_6581 <= 1'h0;
      p2_bit_slice_6582 <= 1'h0;
      p2_bit_slice_6583 <= 1'h0;
      p2_bit_slice_6584 <= 1'h0;
      p2_bit_slice_6585 <= 1'h0;
      p2_bit_slice_6586 <= 1'h0;
      p2_bit_slice_6587 <= 1'h0;
      p2_bit_slice_6588 <= 1'h0;
      p2_bit_slice_6589 <= 1'h0;
      p2_bit_slice_6590 <= 1'h0;
      p2_bit_slice_6591 <= 1'h0;
      p2_bit_slice_6592 <= 1'h0;
      p2_bit_slice_6593 <= 1'h0;
      p2_bit_slice_6594 <= 1'h0;
      p2_bit_slice_6595 <= 1'h0;
      p2_bit_slice_6596 <= 1'h0;
      p2_bit_slice_6597 <= 1'h0;
      p2_bit_slice_6598 <= 1'h0;
      p2_bit_slice_6599 <= 1'h0;
      p2_bit_slice_6600 <= 1'h0;
      p2_bit_slice_6601 <= 1'h0;
      p2_bit_slice_6602 <= 1'h0;
      p2_bit_slice_6603 <= 1'h0;
      p2_bit_slice_6604 <= 1'h0;
      p2_bit_slice_6605 <= 1'h0;
      p2_bit_slice_6606 <= 1'h0;
      p2_bit_slice_6607 <= 1'h0;
      p2_negated <= 1'h0;
      p3_b <= 32'h0000_0000;
      p3_uge_6683 <= 1'h0;
      p3_bivisor__1 <= 33'h0_0000_0000;
      p3_uge_6691 <= 1'h0;
      p3_uge_6771 <= 1'h0;
      p3_concat_6850 <= 32'h0000_0000;
      p3_uge_6851 <= 1'h0;
      p3_bit_slice_6580 <= 1'h0;
      p3_bit_slice_6581 <= 1'h0;
      p3_bit_slice_6582 <= 1'h0;
      p3_bit_slice_6583 <= 1'h0;
      p3_bit_slice_6584 <= 1'h0;
      p3_bit_slice_6585 <= 1'h0;
      p3_bit_slice_6586 <= 1'h0;
      p3_bit_slice_6587 <= 1'h0;
      p3_bit_slice_6588 <= 1'h0;
      p3_bit_slice_6589 <= 1'h0;
      p3_bit_slice_6590 <= 1'h0;
      p3_bit_slice_6591 <= 1'h0;
      p3_bit_slice_6592 <= 1'h0;
      p3_bit_slice_6593 <= 1'h0;
      p3_bit_slice_6594 <= 1'h0;
      p3_bit_slice_6595 <= 1'h0;
      p3_bit_slice_6596 <= 1'h0;
      p3_bit_slice_6597 <= 1'h0;
      p3_bit_slice_6598 <= 1'h0;
      p3_bit_slice_6599 <= 1'h0;
      p3_bit_slice_6600 <= 1'h0;
      p3_bit_slice_6601 <= 1'h0;
      p3_bit_slice_6602 <= 1'h0;
      p3_bit_slice_6603 <= 1'h0;
      p3_bit_slice_6604 <= 1'h0;
      p3_bit_slice_6605 <= 1'h0;
      p3_bit_slice_6606 <= 1'h0;
      p3_bit_slice_6607 <= 1'h0;
      p3_negated <= 1'h0;
      p4_b <= 32'h0000_0000;
      p4_uge_6683 <= 1'h0;
      p4_bivisor__1 <= 33'h0_0000_0000;
      p4_uge_6691 <= 1'h0;
      p4_uge_6771 <= 1'h0;
      p4_uge_6851 <= 1'h0;
      p4_concat_6930 <= 32'h0000_0000;
      p4_uge_6931 <= 1'h0;
      p4_bit_slice_6581 <= 1'h0;
      p4_bit_slice_6582 <= 1'h0;
      p4_bit_slice_6583 <= 1'h0;
      p4_bit_slice_6584 <= 1'h0;
      p4_bit_slice_6585 <= 1'h0;
      p4_bit_slice_6586 <= 1'h0;
      p4_bit_slice_6587 <= 1'h0;
      p4_bit_slice_6588 <= 1'h0;
      p4_bit_slice_6589 <= 1'h0;
      p4_bit_slice_6590 <= 1'h0;
      p4_bit_slice_6591 <= 1'h0;
      p4_bit_slice_6592 <= 1'h0;
      p4_bit_slice_6593 <= 1'h0;
      p4_bit_slice_6594 <= 1'h0;
      p4_bit_slice_6595 <= 1'h0;
      p4_bit_slice_6596 <= 1'h0;
      p4_bit_slice_6597 <= 1'h0;
      p4_bit_slice_6598 <= 1'h0;
      p4_bit_slice_6599 <= 1'h0;
      p4_bit_slice_6600 <= 1'h0;
      p4_bit_slice_6601 <= 1'h0;
      p4_bit_slice_6602 <= 1'h0;
      p4_bit_slice_6603 <= 1'h0;
      p4_bit_slice_6604 <= 1'h0;
      p4_bit_slice_6605 <= 1'h0;
      p4_bit_slice_6606 <= 1'h0;
      p4_bit_slice_6607 <= 1'h0;
      p4_negated <= 1'h0;
      p5_b <= 32'h0000_0000;
      p5_uge_6683 <= 1'h0;
      p5_bivisor__1 <= 33'h0_0000_0000;
      p5_uge_6691 <= 1'h0;
      p5_uge_6771 <= 1'h0;
      p5_uge_6851 <= 1'h0;
      p5_uge_6931 <= 1'h0;
      p5_concat_7010 <= 32'h0000_0000;
      p5_uge_7011 <= 1'h0;
      p5_bit_slice_6582 <= 1'h0;
      p5_bit_slice_6583 <= 1'h0;
      p5_bit_slice_6584 <= 1'h0;
      p5_bit_slice_6585 <= 1'h0;
      p5_bit_slice_6586 <= 1'h0;
      p5_bit_slice_6587 <= 1'h0;
      p5_bit_slice_6588 <= 1'h0;
      p5_bit_slice_6589 <= 1'h0;
      p5_bit_slice_6590 <= 1'h0;
      p5_bit_slice_6591 <= 1'h0;
      p5_bit_slice_6592 <= 1'h0;
      p5_bit_slice_6593 <= 1'h0;
      p5_bit_slice_6594 <= 1'h0;
      p5_bit_slice_6595 <= 1'h0;
      p5_bit_slice_6596 <= 1'h0;
      p5_bit_slice_6597 <= 1'h0;
      p5_bit_slice_6598 <= 1'h0;
      p5_bit_slice_6599 <= 1'h0;
      p5_bit_slice_6600 <= 1'h0;
      p5_bit_slice_6601 <= 1'h0;
      p5_bit_slice_6602 <= 1'h0;
      p5_bit_slice_6603 <= 1'h0;
      p5_bit_slice_6604 <= 1'h0;
      p5_bit_slice_6605 <= 1'h0;
      p5_bit_slice_6606 <= 1'h0;
      p5_bit_slice_6607 <= 1'h0;
      p5_negated <= 1'h0;
      p6_b <= 32'h0000_0000;
      p6_uge_6683 <= 1'h0;
      p6_bivisor__1 <= 33'h0_0000_0000;
      p6_uge_6691 <= 1'h0;
      p6_uge_6771 <= 1'h0;
      p6_uge_6851 <= 1'h0;
      p6_uge_6931 <= 1'h0;
      p6_uge_7011 <= 1'h0;
      p6_concat_7090 <= 32'h0000_0000;
      p6_uge_7091 <= 1'h0;
      p6_bit_slice_6583 <= 1'h0;
      p6_bit_slice_6584 <= 1'h0;
      p6_bit_slice_6585 <= 1'h0;
      p6_bit_slice_6586 <= 1'h0;
      p6_bit_slice_6587 <= 1'h0;
      p6_bit_slice_6588 <= 1'h0;
      p6_bit_slice_6589 <= 1'h0;
      p6_bit_slice_6590 <= 1'h0;
      p6_bit_slice_6591 <= 1'h0;
      p6_bit_slice_6592 <= 1'h0;
      p6_bit_slice_6593 <= 1'h0;
      p6_bit_slice_6594 <= 1'h0;
      p6_bit_slice_6595 <= 1'h0;
      p6_bit_slice_6596 <= 1'h0;
      p6_bit_slice_6597 <= 1'h0;
      p6_bit_slice_6598 <= 1'h0;
      p6_bit_slice_6599 <= 1'h0;
      p6_bit_slice_6600 <= 1'h0;
      p6_bit_slice_6601 <= 1'h0;
      p6_bit_slice_6602 <= 1'h0;
      p6_bit_slice_6603 <= 1'h0;
      p6_bit_slice_6604 <= 1'h0;
      p6_bit_slice_6605 <= 1'h0;
      p6_bit_slice_6606 <= 1'h0;
      p6_bit_slice_6607 <= 1'h0;
      p6_negated <= 1'h0;
      p7_b <= 32'h0000_0000;
      p7_uge_6683 <= 1'h0;
      p7_bivisor__1 <= 33'h0_0000_0000;
      p7_uge_6691 <= 1'h0;
      p7_uge_6771 <= 1'h0;
      p7_uge_6851 <= 1'h0;
      p7_uge_6931 <= 1'h0;
      p7_uge_7011 <= 1'h0;
      p7_uge_7091 <= 1'h0;
      p7_concat_7170 <= 32'h0000_0000;
      p7_uge_7171 <= 1'h0;
      p7_bit_slice_6584 <= 1'h0;
      p7_bit_slice_6585 <= 1'h0;
      p7_bit_slice_6586 <= 1'h0;
      p7_bit_slice_6587 <= 1'h0;
      p7_bit_slice_6588 <= 1'h0;
      p7_bit_slice_6589 <= 1'h0;
      p7_bit_slice_6590 <= 1'h0;
      p7_bit_slice_6591 <= 1'h0;
      p7_bit_slice_6592 <= 1'h0;
      p7_bit_slice_6593 <= 1'h0;
      p7_bit_slice_6594 <= 1'h0;
      p7_bit_slice_6595 <= 1'h0;
      p7_bit_slice_6596 <= 1'h0;
      p7_bit_slice_6597 <= 1'h0;
      p7_bit_slice_6598 <= 1'h0;
      p7_bit_slice_6599 <= 1'h0;
      p7_bit_slice_6600 <= 1'h0;
      p7_bit_slice_6601 <= 1'h0;
      p7_bit_slice_6602 <= 1'h0;
      p7_bit_slice_6603 <= 1'h0;
      p7_bit_slice_6604 <= 1'h0;
      p7_bit_slice_6605 <= 1'h0;
      p7_bit_slice_6606 <= 1'h0;
      p7_bit_slice_6607 <= 1'h0;
      p7_negated <= 1'h0;
      p8_b <= 32'h0000_0000;
      p8_uge_6683 <= 1'h0;
      p8_bivisor__1 <= 33'h0_0000_0000;
      p8_uge_6691 <= 1'h0;
      p8_uge_6771 <= 1'h0;
      p8_uge_6851 <= 1'h0;
      p8_uge_6931 <= 1'h0;
      p8_uge_7011 <= 1'h0;
      p8_uge_7091 <= 1'h0;
      p8_uge_7171 <= 1'h0;
      p8_concat_7250 <= 32'h0000_0000;
      p8_uge_7251 <= 1'h0;
      p8_bit_slice_6585 <= 1'h0;
      p8_bit_slice_6586 <= 1'h0;
      p8_bit_slice_6587 <= 1'h0;
      p8_bit_slice_6588 <= 1'h0;
      p8_bit_slice_6589 <= 1'h0;
      p8_bit_slice_6590 <= 1'h0;
      p8_bit_slice_6591 <= 1'h0;
      p8_bit_slice_6592 <= 1'h0;
      p8_bit_slice_6593 <= 1'h0;
      p8_bit_slice_6594 <= 1'h0;
      p8_bit_slice_6595 <= 1'h0;
      p8_bit_slice_6596 <= 1'h0;
      p8_bit_slice_6597 <= 1'h0;
      p8_bit_slice_6598 <= 1'h0;
      p8_bit_slice_6599 <= 1'h0;
      p8_bit_slice_6600 <= 1'h0;
      p8_bit_slice_6601 <= 1'h0;
      p8_bit_slice_6602 <= 1'h0;
      p8_bit_slice_6603 <= 1'h0;
      p8_bit_slice_6604 <= 1'h0;
      p8_bit_slice_6605 <= 1'h0;
      p8_bit_slice_6606 <= 1'h0;
      p8_bit_slice_6607 <= 1'h0;
      p8_negated <= 1'h0;
      p9_b <= 32'h0000_0000;
      p9_uge_6683 <= 1'h0;
      p9_bivisor__1 <= 33'h0_0000_0000;
      p9_uge_6691 <= 1'h0;
      p9_uge_6771 <= 1'h0;
      p9_uge_6851 <= 1'h0;
      p9_uge_6931 <= 1'h0;
      p9_uge_7011 <= 1'h0;
      p9_uge_7091 <= 1'h0;
      p9_uge_7171 <= 1'h0;
      p9_uge_7251 <= 1'h0;
      p9_concat_7330 <= 32'h0000_0000;
      p9_uge_7331 <= 1'h0;
      p9_bit_slice_6586 <= 1'h0;
      p9_bit_slice_6587 <= 1'h0;
      p9_bit_slice_6588 <= 1'h0;
      p9_bit_slice_6589 <= 1'h0;
      p9_bit_slice_6590 <= 1'h0;
      p9_bit_slice_6591 <= 1'h0;
      p9_bit_slice_6592 <= 1'h0;
      p9_bit_slice_6593 <= 1'h0;
      p9_bit_slice_6594 <= 1'h0;
      p9_bit_slice_6595 <= 1'h0;
      p9_bit_slice_6596 <= 1'h0;
      p9_bit_slice_6597 <= 1'h0;
      p9_bit_slice_6598 <= 1'h0;
      p9_bit_slice_6599 <= 1'h0;
      p9_bit_slice_6600 <= 1'h0;
      p9_bit_slice_6601 <= 1'h0;
      p9_bit_slice_6602 <= 1'h0;
      p9_bit_slice_6603 <= 1'h0;
      p9_bit_slice_6604 <= 1'h0;
      p9_bit_slice_6605 <= 1'h0;
      p9_bit_slice_6606 <= 1'h0;
      p9_bit_slice_6607 <= 1'h0;
      p9_negated <= 1'h0;
      p10_b <= 32'h0000_0000;
      p10_uge_6683 <= 1'h0;
      p10_bivisor__1 <= 33'h0_0000_0000;
      p10_uge_6691 <= 1'h0;
      p10_uge_6771 <= 1'h0;
      p10_uge_6851 <= 1'h0;
      p10_uge_6931 <= 1'h0;
      p10_uge_7011 <= 1'h0;
      p10_uge_7091 <= 1'h0;
      p10_uge_7171 <= 1'h0;
      p10_uge_7251 <= 1'h0;
      p10_uge_7331 <= 1'h0;
      p10_concat_7410 <= 32'h0000_0000;
      p10_uge_7411 <= 1'h0;
      p10_bit_slice_6587 <= 1'h0;
      p10_bit_slice_6588 <= 1'h0;
      p10_bit_slice_6589 <= 1'h0;
      p10_bit_slice_6590 <= 1'h0;
      p10_bit_slice_6591 <= 1'h0;
      p10_bit_slice_6592 <= 1'h0;
      p10_bit_slice_6593 <= 1'h0;
      p10_bit_slice_6594 <= 1'h0;
      p10_bit_slice_6595 <= 1'h0;
      p10_bit_slice_6596 <= 1'h0;
      p10_bit_slice_6597 <= 1'h0;
      p10_bit_slice_6598 <= 1'h0;
      p10_bit_slice_6599 <= 1'h0;
      p10_bit_slice_6600 <= 1'h0;
      p10_bit_slice_6601 <= 1'h0;
      p10_bit_slice_6602 <= 1'h0;
      p10_bit_slice_6603 <= 1'h0;
      p10_bit_slice_6604 <= 1'h0;
      p10_bit_slice_6605 <= 1'h0;
      p10_bit_slice_6606 <= 1'h0;
      p10_bit_slice_6607 <= 1'h0;
      p10_negated <= 1'h0;
      p11_b <= 32'h0000_0000;
      p11_uge_6683 <= 1'h0;
      p11_bivisor__1 <= 33'h0_0000_0000;
      p11_uge_6691 <= 1'h0;
      p11_uge_6771 <= 1'h0;
      p11_uge_6851 <= 1'h0;
      p11_uge_6931 <= 1'h0;
      p11_uge_7011 <= 1'h0;
      p11_uge_7091 <= 1'h0;
      p11_uge_7171 <= 1'h0;
      p11_uge_7251 <= 1'h0;
      p11_uge_7331 <= 1'h0;
      p11_uge_7411 <= 1'h0;
      p11_concat_7490 <= 32'h0000_0000;
      p11_uge_7491 <= 1'h0;
      p11_bit_slice_6588 <= 1'h0;
      p11_bit_slice_6589 <= 1'h0;
      p11_bit_slice_6590 <= 1'h0;
      p11_bit_slice_6591 <= 1'h0;
      p11_bit_slice_6592 <= 1'h0;
      p11_bit_slice_6593 <= 1'h0;
      p11_bit_slice_6594 <= 1'h0;
      p11_bit_slice_6595 <= 1'h0;
      p11_bit_slice_6596 <= 1'h0;
      p11_bit_slice_6597 <= 1'h0;
      p11_bit_slice_6598 <= 1'h0;
      p11_bit_slice_6599 <= 1'h0;
      p11_bit_slice_6600 <= 1'h0;
      p11_bit_slice_6601 <= 1'h0;
      p11_bit_slice_6602 <= 1'h0;
      p11_bit_slice_6603 <= 1'h0;
      p11_bit_slice_6604 <= 1'h0;
      p11_bit_slice_6605 <= 1'h0;
      p11_bit_slice_6606 <= 1'h0;
      p11_bit_slice_6607 <= 1'h0;
      p11_negated <= 1'h0;
      p12_b <= 32'h0000_0000;
      p12_uge_6683 <= 1'h0;
      p12_bivisor__1 <= 33'h0_0000_0000;
      p12_uge_6691 <= 1'h0;
      p12_uge_6771 <= 1'h0;
      p12_uge_6851 <= 1'h0;
      p12_uge_6931 <= 1'h0;
      p12_uge_7011 <= 1'h0;
      p12_uge_7091 <= 1'h0;
      p12_uge_7171 <= 1'h0;
      p12_uge_7251 <= 1'h0;
      p12_uge_7331 <= 1'h0;
      p12_uge_7411 <= 1'h0;
      p12_uge_7491 <= 1'h0;
      p12_concat_7570 <= 32'h0000_0000;
      p12_uge_7571 <= 1'h0;
      p12_bit_slice_6589 <= 1'h0;
      p12_bit_slice_6590 <= 1'h0;
      p12_bit_slice_6591 <= 1'h0;
      p12_bit_slice_6592 <= 1'h0;
      p12_bit_slice_6593 <= 1'h0;
      p12_bit_slice_6594 <= 1'h0;
      p12_bit_slice_6595 <= 1'h0;
      p12_bit_slice_6596 <= 1'h0;
      p12_bit_slice_6597 <= 1'h0;
      p12_bit_slice_6598 <= 1'h0;
      p12_bit_slice_6599 <= 1'h0;
      p12_bit_slice_6600 <= 1'h0;
      p12_bit_slice_6601 <= 1'h0;
      p12_bit_slice_6602 <= 1'h0;
      p12_bit_slice_6603 <= 1'h0;
      p12_bit_slice_6604 <= 1'h0;
      p12_bit_slice_6605 <= 1'h0;
      p12_bit_slice_6606 <= 1'h0;
      p12_bit_slice_6607 <= 1'h0;
      p12_negated <= 1'h0;
      p13_b <= 32'h0000_0000;
      p13_uge_6683 <= 1'h0;
      p13_bivisor__1 <= 33'h0_0000_0000;
      p13_uge_6691 <= 1'h0;
      p13_uge_6771 <= 1'h0;
      p13_uge_6851 <= 1'h0;
      p13_uge_6931 <= 1'h0;
      p13_uge_7011 <= 1'h0;
      p13_uge_7091 <= 1'h0;
      p13_uge_7171 <= 1'h0;
      p13_uge_7251 <= 1'h0;
      p13_uge_7331 <= 1'h0;
      p13_uge_7411 <= 1'h0;
      p13_uge_7491 <= 1'h0;
      p13_uge_7571 <= 1'h0;
      p13_concat_7650 <= 32'h0000_0000;
      p13_uge_7651 <= 1'h0;
      p13_bit_slice_6590 <= 1'h0;
      p13_bit_slice_6591 <= 1'h0;
      p13_bit_slice_6592 <= 1'h0;
      p13_bit_slice_6593 <= 1'h0;
      p13_bit_slice_6594 <= 1'h0;
      p13_bit_slice_6595 <= 1'h0;
      p13_bit_slice_6596 <= 1'h0;
      p13_bit_slice_6597 <= 1'h0;
      p13_bit_slice_6598 <= 1'h0;
      p13_bit_slice_6599 <= 1'h0;
      p13_bit_slice_6600 <= 1'h0;
      p13_bit_slice_6601 <= 1'h0;
      p13_bit_slice_6602 <= 1'h0;
      p13_bit_slice_6603 <= 1'h0;
      p13_bit_slice_6604 <= 1'h0;
      p13_bit_slice_6605 <= 1'h0;
      p13_bit_slice_6606 <= 1'h0;
      p13_bit_slice_6607 <= 1'h0;
      p13_negated <= 1'h0;
      p14_b <= 32'h0000_0000;
      p14_uge_6683 <= 1'h0;
      p14_bivisor__1 <= 33'h0_0000_0000;
      p14_uge_6691 <= 1'h0;
      p14_uge_6771 <= 1'h0;
      p14_uge_6851 <= 1'h0;
      p14_uge_6931 <= 1'h0;
      p14_uge_7011 <= 1'h0;
      p14_uge_7091 <= 1'h0;
      p14_uge_7171 <= 1'h0;
      p14_uge_7251 <= 1'h0;
      p14_uge_7331 <= 1'h0;
      p14_uge_7411 <= 1'h0;
      p14_uge_7491 <= 1'h0;
      p14_uge_7571 <= 1'h0;
      p14_uge_7651 <= 1'h0;
      p14_concat_7730 <= 32'h0000_0000;
      p14_uge_7731 <= 1'h0;
      p14_bit_slice_6591 <= 1'h0;
      p14_bit_slice_6592 <= 1'h0;
      p14_bit_slice_6593 <= 1'h0;
      p14_bit_slice_6594 <= 1'h0;
      p14_bit_slice_6595 <= 1'h0;
      p14_bit_slice_6596 <= 1'h0;
      p14_bit_slice_6597 <= 1'h0;
      p14_bit_slice_6598 <= 1'h0;
      p14_bit_slice_6599 <= 1'h0;
      p14_bit_slice_6600 <= 1'h0;
      p14_bit_slice_6601 <= 1'h0;
      p14_bit_slice_6602 <= 1'h0;
      p14_bit_slice_6603 <= 1'h0;
      p14_bit_slice_6604 <= 1'h0;
      p14_bit_slice_6605 <= 1'h0;
      p14_bit_slice_6606 <= 1'h0;
      p14_bit_slice_6607 <= 1'h0;
      p14_negated <= 1'h0;
      p15_b <= 32'h0000_0000;
      p15_uge_6683 <= 1'h0;
      p15_bivisor__1 <= 33'h0_0000_0000;
      p15_uge_6691 <= 1'h0;
      p15_uge_6771 <= 1'h0;
      p15_uge_6851 <= 1'h0;
      p15_uge_6931 <= 1'h0;
      p15_uge_7011 <= 1'h0;
      p15_uge_7091 <= 1'h0;
      p15_uge_7171 <= 1'h0;
      p15_uge_7251 <= 1'h0;
      p15_uge_7331 <= 1'h0;
      p15_uge_7411 <= 1'h0;
      p15_uge_7491 <= 1'h0;
      p15_uge_7571 <= 1'h0;
      p15_uge_7651 <= 1'h0;
      p15_uge_7731 <= 1'h0;
      p15_concat_7810 <= 32'h0000_0000;
      p15_uge_7811 <= 1'h0;
      p15_bit_slice_6592 <= 1'h0;
      p15_bit_slice_6593 <= 1'h0;
      p15_bit_slice_6594 <= 1'h0;
      p15_bit_slice_6595 <= 1'h0;
      p15_bit_slice_6596 <= 1'h0;
      p15_bit_slice_6597 <= 1'h0;
      p15_bit_slice_6598 <= 1'h0;
      p15_bit_slice_6599 <= 1'h0;
      p15_bit_slice_6600 <= 1'h0;
      p15_bit_slice_6601 <= 1'h0;
      p15_bit_slice_6602 <= 1'h0;
      p15_bit_slice_6603 <= 1'h0;
      p15_bit_slice_6604 <= 1'h0;
      p15_bit_slice_6605 <= 1'h0;
      p15_bit_slice_6606 <= 1'h0;
      p15_bit_slice_6607 <= 1'h0;
      p15_negated <= 1'h0;
      p16_b <= 32'h0000_0000;
      p16_uge_6683 <= 1'h0;
      p16_bivisor__1 <= 33'h0_0000_0000;
      p16_uge_6691 <= 1'h0;
      p16_uge_6771 <= 1'h0;
      p16_uge_6851 <= 1'h0;
      p16_uge_6931 <= 1'h0;
      p16_uge_7011 <= 1'h0;
      p16_uge_7091 <= 1'h0;
      p16_uge_7171 <= 1'h0;
      p16_uge_7251 <= 1'h0;
      p16_uge_7331 <= 1'h0;
      p16_uge_7411 <= 1'h0;
      p16_uge_7491 <= 1'h0;
      p16_uge_7571 <= 1'h0;
      p16_uge_7651 <= 1'h0;
      p16_uge_7731 <= 1'h0;
      p16_uge_7811 <= 1'h0;
      p16_concat_7890 <= 32'h0000_0000;
      p16_uge_7891 <= 1'h0;
      p16_bit_slice_6593 <= 1'h0;
      p16_bit_slice_6594 <= 1'h0;
      p16_bit_slice_6595 <= 1'h0;
      p16_bit_slice_6596 <= 1'h0;
      p16_bit_slice_6597 <= 1'h0;
      p16_bit_slice_6598 <= 1'h0;
      p16_bit_slice_6599 <= 1'h0;
      p16_bit_slice_6600 <= 1'h0;
      p16_bit_slice_6601 <= 1'h0;
      p16_bit_slice_6602 <= 1'h0;
      p16_bit_slice_6603 <= 1'h0;
      p16_bit_slice_6604 <= 1'h0;
      p16_bit_slice_6605 <= 1'h0;
      p16_bit_slice_6606 <= 1'h0;
      p16_bit_slice_6607 <= 1'h0;
      p16_negated <= 1'h0;
      p17_b <= 32'h0000_0000;
      p17_uge_6683 <= 1'h0;
      p17_bivisor__1 <= 33'h0_0000_0000;
      p17_uge_6691 <= 1'h0;
      p17_uge_6771 <= 1'h0;
      p17_uge_6851 <= 1'h0;
      p17_uge_6931 <= 1'h0;
      p17_uge_7011 <= 1'h0;
      p17_uge_7091 <= 1'h0;
      p17_uge_7171 <= 1'h0;
      p17_uge_7251 <= 1'h0;
      p17_uge_7331 <= 1'h0;
      p17_uge_7411 <= 1'h0;
      p17_uge_7491 <= 1'h0;
      p17_uge_7571 <= 1'h0;
      p17_uge_7651 <= 1'h0;
      p17_uge_7731 <= 1'h0;
      p17_uge_7811 <= 1'h0;
      p17_uge_7891 <= 1'h0;
      p17_concat_7970 <= 32'h0000_0000;
      p17_uge_7971 <= 1'h0;
      p17_bit_slice_6594 <= 1'h0;
      p17_bit_slice_6595 <= 1'h0;
      p17_bit_slice_6596 <= 1'h0;
      p17_bit_slice_6597 <= 1'h0;
      p17_bit_slice_6598 <= 1'h0;
      p17_bit_slice_6599 <= 1'h0;
      p17_bit_slice_6600 <= 1'h0;
      p17_bit_slice_6601 <= 1'h0;
      p17_bit_slice_6602 <= 1'h0;
      p17_bit_slice_6603 <= 1'h0;
      p17_bit_slice_6604 <= 1'h0;
      p17_bit_slice_6605 <= 1'h0;
      p17_bit_slice_6606 <= 1'h0;
      p17_bit_slice_6607 <= 1'h0;
      p17_negated <= 1'h0;
      p18_b <= 32'h0000_0000;
      p18_uge_6683 <= 1'h0;
      p18_bivisor__1 <= 33'h0_0000_0000;
      p18_uge_6691 <= 1'h0;
      p18_uge_6771 <= 1'h0;
      p18_uge_6851 <= 1'h0;
      p18_uge_6931 <= 1'h0;
      p18_uge_7011 <= 1'h0;
      p18_uge_7091 <= 1'h0;
      p18_uge_7171 <= 1'h0;
      p18_uge_7251 <= 1'h0;
      p18_uge_7331 <= 1'h0;
      p18_uge_7411 <= 1'h0;
      p18_uge_7491 <= 1'h0;
      p18_uge_7571 <= 1'h0;
      p18_uge_7651 <= 1'h0;
      p18_uge_7731 <= 1'h0;
      p18_uge_7811 <= 1'h0;
      p18_uge_7891 <= 1'h0;
      p18_uge_7971 <= 1'h0;
      p18_concat_8050 <= 32'h0000_0000;
      p18_uge_8051 <= 1'h0;
      p18_bit_slice_6595 <= 1'h0;
      p18_bit_slice_6596 <= 1'h0;
      p18_bit_slice_6597 <= 1'h0;
      p18_bit_slice_6598 <= 1'h0;
      p18_bit_slice_6599 <= 1'h0;
      p18_bit_slice_6600 <= 1'h0;
      p18_bit_slice_6601 <= 1'h0;
      p18_bit_slice_6602 <= 1'h0;
      p18_bit_slice_6603 <= 1'h0;
      p18_bit_slice_6604 <= 1'h0;
      p18_bit_slice_6605 <= 1'h0;
      p18_bit_slice_6606 <= 1'h0;
      p18_bit_slice_6607 <= 1'h0;
      p18_negated <= 1'h0;
      p19_b <= 32'h0000_0000;
      p19_uge_6683 <= 1'h0;
      p19_bivisor__1 <= 33'h0_0000_0000;
      p19_uge_6691 <= 1'h0;
      p19_uge_6771 <= 1'h0;
      p19_uge_6851 <= 1'h0;
      p19_uge_6931 <= 1'h0;
      p19_uge_7011 <= 1'h0;
      p19_uge_7091 <= 1'h0;
      p19_uge_7171 <= 1'h0;
      p19_uge_7251 <= 1'h0;
      p19_uge_7331 <= 1'h0;
      p19_uge_7411 <= 1'h0;
      p19_uge_7491 <= 1'h0;
      p19_uge_7571 <= 1'h0;
      p19_uge_7651 <= 1'h0;
      p19_uge_7731 <= 1'h0;
      p19_uge_7811 <= 1'h0;
      p19_uge_7891 <= 1'h0;
      p19_uge_7971 <= 1'h0;
      p19_uge_8051 <= 1'h0;
      p19_concat_8130 <= 32'h0000_0000;
      p19_uge_8131 <= 1'h0;
      p19_bit_slice_6596 <= 1'h0;
      p19_bit_slice_6597 <= 1'h0;
      p19_bit_slice_6598 <= 1'h0;
      p19_bit_slice_6599 <= 1'h0;
      p19_bit_slice_6600 <= 1'h0;
      p19_bit_slice_6601 <= 1'h0;
      p19_bit_slice_6602 <= 1'h0;
      p19_bit_slice_6603 <= 1'h0;
      p19_bit_slice_6604 <= 1'h0;
      p19_bit_slice_6605 <= 1'h0;
      p19_bit_slice_6606 <= 1'h0;
      p19_bit_slice_6607 <= 1'h0;
      p19_negated <= 1'h0;
      p20_b <= 32'h0000_0000;
      p20_uge_6683 <= 1'h0;
      p20_bivisor__1 <= 33'h0_0000_0000;
      p20_uge_6691 <= 1'h0;
      p20_uge_6771 <= 1'h0;
      p20_uge_6851 <= 1'h0;
      p20_uge_6931 <= 1'h0;
      p20_uge_7011 <= 1'h0;
      p20_uge_7091 <= 1'h0;
      p20_uge_7171 <= 1'h0;
      p20_uge_7251 <= 1'h0;
      p20_uge_7331 <= 1'h0;
      p20_uge_7411 <= 1'h0;
      p20_uge_7491 <= 1'h0;
      p20_uge_7571 <= 1'h0;
      p20_uge_7651 <= 1'h0;
      p20_uge_7731 <= 1'h0;
      p20_uge_7811 <= 1'h0;
      p20_uge_7891 <= 1'h0;
      p20_uge_7971 <= 1'h0;
      p20_uge_8051 <= 1'h0;
      p20_uge_8131 <= 1'h0;
      p20_concat_8210 <= 32'h0000_0000;
      p20_uge_8211 <= 1'h0;
      p20_bit_slice_6597 <= 1'h0;
      p20_bit_slice_6598 <= 1'h0;
      p20_bit_slice_6599 <= 1'h0;
      p20_bit_slice_6600 <= 1'h0;
      p20_bit_slice_6601 <= 1'h0;
      p20_bit_slice_6602 <= 1'h0;
      p20_bit_slice_6603 <= 1'h0;
      p20_bit_slice_6604 <= 1'h0;
      p20_bit_slice_6605 <= 1'h0;
      p20_bit_slice_6606 <= 1'h0;
      p20_bit_slice_6607 <= 1'h0;
      p20_negated <= 1'h0;
      p21_b <= 32'h0000_0000;
      p21_uge_6683 <= 1'h0;
      p21_bivisor__1 <= 33'h0_0000_0000;
      p21_uge_6691 <= 1'h0;
      p21_uge_6771 <= 1'h0;
      p21_uge_6851 <= 1'h0;
      p21_uge_6931 <= 1'h0;
      p21_uge_7011 <= 1'h0;
      p21_uge_7091 <= 1'h0;
      p21_uge_7171 <= 1'h0;
      p21_uge_7251 <= 1'h0;
      p21_uge_7331 <= 1'h0;
      p21_uge_7411 <= 1'h0;
      p21_uge_7491 <= 1'h0;
      p21_uge_7571 <= 1'h0;
      p21_uge_7651 <= 1'h0;
      p21_uge_7731 <= 1'h0;
      p21_uge_7811 <= 1'h0;
      p21_uge_7891 <= 1'h0;
      p21_uge_7971 <= 1'h0;
      p21_uge_8051 <= 1'h0;
      p21_uge_8131 <= 1'h0;
      p21_uge_8211 <= 1'h0;
      p21_concat_8290 <= 32'h0000_0000;
      p21_uge_8291 <= 1'h0;
      p21_bit_slice_6598 <= 1'h0;
      p21_bit_slice_6599 <= 1'h0;
      p21_bit_slice_6600 <= 1'h0;
      p21_bit_slice_6601 <= 1'h0;
      p21_bit_slice_6602 <= 1'h0;
      p21_bit_slice_6603 <= 1'h0;
      p21_bit_slice_6604 <= 1'h0;
      p21_bit_slice_6605 <= 1'h0;
      p21_bit_slice_6606 <= 1'h0;
      p21_bit_slice_6607 <= 1'h0;
      p21_negated <= 1'h0;
      p22_b <= 32'h0000_0000;
      p22_uge_6683 <= 1'h0;
      p22_bivisor__1 <= 33'h0_0000_0000;
      p22_uge_6691 <= 1'h0;
      p22_uge_6771 <= 1'h0;
      p22_uge_6851 <= 1'h0;
      p22_uge_6931 <= 1'h0;
      p22_uge_7011 <= 1'h0;
      p22_uge_7091 <= 1'h0;
      p22_uge_7171 <= 1'h0;
      p22_uge_7251 <= 1'h0;
      p22_uge_7331 <= 1'h0;
      p22_uge_7411 <= 1'h0;
      p22_uge_7491 <= 1'h0;
      p22_uge_7571 <= 1'h0;
      p22_uge_7651 <= 1'h0;
      p22_uge_7731 <= 1'h0;
      p22_uge_7811 <= 1'h0;
      p22_uge_7891 <= 1'h0;
      p22_uge_7971 <= 1'h0;
      p22_uge_8051 <= 1'h0;
      p22_uge_8131 <= 1'h0;
      p22_uge_8211 <= 1'h0;
      p22_uge_8291 <= 1'h0;
      p22_concat_8370 <= 32'h0000_0000;
      p22_uge_8371 <= 1'h0;
      p22_bit_slice_6599 <= 1'h0;
      p22_bit_slice_6600 <= 1'h0;
      p22_bit_slice_6601 <= 1'h0;
      p22_bit_slice_6602 <= 1'h0;
      p22_bit_slice_6603 <= 1'h0;
      p22_bit_slice_6604 <= 1'h0;
      p22_bit_slice_6605 <= 1'h0;
      p22_bit_slice_6606 <= 1'h0;
      p22_bit_slice_6607 <= 1'h0;
      p22_negated <= 1'h0;
      p23_b <= 32'h0000_0000;
      p23_uge_6683 <= 1'h0;
      p23_bivisor__1 <= 33'h0_0000_0000;
      p23_uge_6691 <= 1'h0;
      p23_uge_6771 <= 1'h0;
      p23_uge_6851 <= 1'h0;
      p23_uge_6931 <= 1'h0;
      p23_uge_7011 <= 1'h0;
      p23_uge_7091 <= 1'h0;
      p23_uge_7171 <= 1'h0;
      p23_uge_7251 <= 1'h0;
      p23_uge_7331 <= 1'h0;
      p23_uge_7411 <= 1'h0;
      p23_uge_7491 <= 1'h0;
      p23_uge_7571 <= 1'h0;
      p23_uge_7651 <= 1'h0;
      p23_uge_7731 <= 1'h0;
      p23_uge_7811 <= 1'h0;
      p23_uge_7891 <= 1'h0;
      p23_uge_7971 <= 1'h0;
      p23_uge_8051 <= 1'h0;
      p23_uge_8131 <= 1'h0;
      p23_uge_8211 <= 1'h0;
      p23_uge_8291 <= 1'h0;
      p23_uge_8371 <= 1'h0;
      p23_concat_8450 <= 32'h0000_0000;
      p23_uge_8451 <= 1'h0;
      p23_bit_slice_6600 <= 1'h0;
      p23_bit_slice_6601 <= 1'h0;
      p23_bit_slice_6602 <= 1'h0;
      p23_bit_slice_6603 <= 1'h0;
      p23_bit_slice_6604 <= 1'h0;
      p23_bit_slice_6605 <= 1'h0;
      p23_bit_slice_6606 <= 1'h0;
      p23_bit_slice_6607 <= 1'h0;
      p23_negated <= 1'h0;
      p24_b <= 32'h0000_0000;
      p24_uge_6683 <= 1'h0;
      p24_bivisor__1 <= 33'h0_0000_0000;
      p24_uge_6691 <= 1'h0;
      p24_uge_6771 <= 1'h0;
      p24_uge_6851 <= 1'h0;
      p24_uge_6931 <= 1'h0;
      p24_uge_7011 <= 1'h0;
      p24_uge_7091 <= 1'h0;
      p24_uge_7171 <= 1'h0;
      p24_uge_7251 <= 1'h0;
      p24_uge_7331 <= 1'h0;
      p24_uge_7411 <= 1'h0;
      p24_uge_7491 <= 1'h0;
      p24_uge_7571 <= 1'h0;
      p24_uge_7651 <= 1'h0;
      p24_uge_7731 <= 1'h0;
      p24_uge_7811 <= 1'h0;
      p24_uge_7891 <= 1'h0;
      p24_uge_7971 <= 1'h0;
      p24_uge_8051 <= 1'h0;
      p24_uge_8131 <= 1'h0;
      p24_uge_8211 <= 1'h0;
      p24_uge_8291 <= 1'h0;
      p24_uge_8371 <= 1'h0;
      p24_uge_8451 <= 1'h0;
      p24_concat_8530 <= 32'h0000_0000;
      p24_uge_8531 <= 1'h0;
      p24_bit_slice_6601 <= 1'h0;
      p24_bit_slice_6602 <= 1'h0;
      p24_bit_slice_6603 <= 1'h0;
      p24_bit_slice_6604 <= 1'h0;
      p24_bit_slice_6605 <= 1'h0;
      p24_bit_slice_6606 <= 1'h0;
      p24_bit_slice_6607 <= 1'h0;
      p24_negated <= 1'h0;
      p25_b <= 32'h0000_0000;
      p25_uge_6683 <= 1'h0;
      p25_bivisor__1 <= 33'h0_0000_0000;
      p25_uge_6691 <= 1'h0;
      p25_uge_6771 <= 1'h0;
      p25_uge_6851 <= 1'h0;
      p25_uge_6931 <= 1'h0;
      p25_uge_7011 <= 1'h0;
      p25_uge_7091 <= 1'h0;
      p25_uge_7171 <= 1'h0;
      p25_uge_7251 <= 1'h0;
      p25_uge_7331 <= 1'h0;
      p25_uge_7411 <= 1'h0;
      p25_uge_7491 <= 1'h0;
      p25_uge_7571 <= 1'h0;
      p25_uge_7651 <= 1'h0;
      p25_uge_7731 <= 1'h0;
      p25_uge_7811 <= 1'h0;
      p25_uge_7891 <= 1'h0;
      p25_uge_7971 <= 1'h0;
      p25_uge_8051 <= 1'h0;
      p25_uge_8131 <= 1'h0;
      p25_uge_8211 <= 1'h0;
      p25_uge_8291 <= 1'h0;
      p25_uge_8371 <= 1'h0;
      p25_uge_8451 <= 1'h0;
      p25_uge_8531 <= 1'h0;
      p25_concat_8610 <= 32'h0000_0000;
      p25_uge_8611 <= 1'h0;
      p25_bit_slice_6602 <= 1'h0;
      p25_bit_slice_6603 <= 1'h0;
      p25_bit_slice_6604 <= 1'h0;
      p25_bit_slice_6605 <= 1'h0;
      p25_bit_slice_6606 <= 1'h0;
      p25_bit_slice_6607 <= 1'h0;
      p25_negated <= 1'h0;
      p26_b <= 32'h0000_0000;
      p26_uge_6683 <= 1'h0;
      p26_bivisor__1 <= 33'h0_0000_0000;
      p26_uge_6691 <= 1'h0;
      p26_uge_6771 <= 1'h0;
      p26_uge_6851 <= 1'h0;
      p26_uge_6931 <= 1'h0;
      p26_uge_7011 <= 1'h0;
      p26_uge_7091 <= 1'h0;
      p26_uge_7171 <= 1'h0;
      p26_uge_7251 <= 1'h0;
      p26_uge_7331 <= 1'h0;
      p26_uge_7411 <= 1'h0;
      p26_uge_7491 <= 1'h0;
      p26_uge_7571 <= 1'h0;
      p26_uge_7651 <= 1'h0;
      p26_uge_7731 <= 1'h0;
      p26_uge_7811 <= 1'h0;
      p26_uge_7891 <= 1'h0;
      p26_uge_7971 <= 1'h0;
      p26_uge_8051 <= 1'h0;
      p26_uge_8131 <= 1'h0;
      p26_uge_8211 <= 1'h0;
      p26_uge_8291 <= 1'h0;
      p26_uge_8371 <= 1'h0;
      p26_uge_8451 <= 1'h0;
      p26_uge_8531 <= 1'h0;
      p26_uge_8611 <= 1'h0;
      p26_concat_8690 <= 32'h0000_0000;
      p26_uge_8691 <= 1'h0;
      p26_bit_slice_6603 <= 1'h0;
      p26_bit_slice_6604 <= 1'h0;
      p26_bit_slice_6605 <= 1'h0;
      p26_bit_slice_6606 <= 1'h0;
      p26_bit_slice_6607 <= 1'h0;
      p26_negated <= 1'h0;
      p27_b <= 32'h0000_0000;
      p27_uge_6683 <= 1'h0;
      p27_bivisor__1 <= 33'h0_0000_0000;
      p27_uge_6691 <= 1'h0;
      p27_uge_6771 <= 1'h0;
      p27_uge_6851 <= 1'h0;
      p27_uge_6931 <= 1'h0;
      p27_uge_7011 <= 1'h0;
      p27_uge_7091 <= 1'h0;
      p27_uge_7171 <= 1'h0;
      p27_uge_7251 <= 1'h0;
      p27_uge_7331 <= 1'h0;
      p27_uge_7411 <= 1'h0;
      p27_uge_7491 <= 1'h0;
      p27_uge_7571 <= 1'h0;
      p27_uge_7651 <= 1'h0;
      p27_uge_7731 <= 1'h0;
      p27_uge_7811 <= 1'h0;
      p27_uge_7891 <= 1'h0;
      p27_uge_7971 <= 1'h0;
      p27_uge_8051 <= 1'h0;
      p27_uge_8131 <= 1'h0;
      p27_uge_8211 <= 1'h0;
      p27_uge_8291 <= 1'h0;
      p27_uge_8371 <= 1'h0;
      p27_uge_8451 <= 1'h0;
      p27_uge_8531 <= 1'h0;
      p27_uge_8611 <= 1'h0;
      p27_uge_8691 <= 1'h0;
      p27_concat_8770 <= 32'h0000_0000;
      p27_uge_8771 <= 1'h0;
      p27_bit_slice_6604 <= 1'h0;
      p27_bit_slice_6605 <= 1'h0;
      p27_bit_slice_6606 <= 1'h0;
      p27_bit_slice_6607 <= 1'h0;
      p27_negated <= 1'h0;
      p28_b <= 32'h0000_0000;
      p28_uge_6683 <= 1'h0;
      p28_bivisor__1 <= 33'h0_0000_0000;
      p28_uge_6691 <= 1'h0;
      p28_uge_6771 <= 1'h0;
      p28_uge_6851 <= 1'h0;
      p28_uge_6931 <= 1'h0;
      p28_uge_7011 <= 1'h0;
      p28_uge_7091 <= 1'h0;
      p28_uge_7171 <= 1'h0;
      p28_uge_7251 <= 1'h0;
      p28_uge_7331 <= 1'h0;
      p28_uge_7411 <= 1'h0;
      p28_uge_7491 <= 1'h0;
      p28_uge_7571 <= 1'h0;
      p28_uge_7651 <= 1'h0;
      p28_uge_7731 <= 1'h0;
      p28_uge_7811 <= 1'h0;
      p28_uge_7891 <= 1'h0;
      p28_uge_7971 <= 1'h0;
      p28_uge_8051 <= 1'h0;
      p28_uge_8131 <= 1'h0;
      p28_uge_8211 <= 1'h0;
      p28_uge_8291 <= 1'h0;
      p28_uge_8371 <= 1'h0;
      p28_uge_8451 <= 1'h0;
      p28_uge_8531 <= 1'h0;
      p28_uge_8611 <= 1'h0;
      p28_uge_8691 <= 1'h0;
      p28_uge_8771 <= 1'h0;
      p28_concat_8850 <= 32'h0000_0000;
      p28_uge_8851 <= 1'h0;
      p28_bit_slice_6605 <= 1'h0;
      p28_bit_slice_6606 <= 1'h0;
      p28_bit_slice_6607 <= 1'h0;
      p28_negated <= 1'h0;
      p29_b <= 32'h0000_0000;
      p29_uge_6683 <= 1'h0;
      p29_bivisor__1 <= 33'h0_0000_0000;
      p29_uge_6691 <= 1'h0;
      p29_uge_6771 <= 1'h0;
      p29_uge_6851 <= 1'h0;
      p29_uge_6931 <= 1'h0;
      p29_uge_7011 <= 1'h0;
      p29_uge_7091 <= 1'h0;
      p29_uge_7171 <= 1'h0;
      p29_uge_7251 <= 1'h0;
      p29_uge_7331 <= 1'h0;
      p29_uge_7411 <= 1'h0;
      p29_uge_7491 <= 1'h0;
      p29_uge_7571 <= 1'h0;
      p29_uge_7651 <= 1'h0;
      p29_uge_7731 <= 1'h0;
      p29_uge_7811 <= 1'h0;
      p29_uge_7891 <= 1'h0;
      p29_uge_7971 <= 1'h0;
      p29_uge_8051 <= 1'h0;
      p29_uge_8131 <= 1'h0;
      p29_uge_8211 <= 1'h0;
      p29_uge_8291 <= 1'h0;
      p29_uge_8371 <= 1'h0;
      p29_uge_8451 <= 1'h0;
      p29_uge_8531 <= 1'h0;
      p29_uge_8611 <= 1'h0;
      p29_uge_8691 <= 1'h0;
      p29_uge_8771 <= 1'h0;
      p29_uge_8851 <= 1'h0;
      p29_concat_8930 <= 32'h0000_0000;
      p29_uge_8931 <= 1'h0;
      p29_bit_slice_6606 <= 1'h0;
      p29_bit_slice_6607 <= 1'h0;
      p29_negated <= 1'h0;
      p30_b <= 32'h0000_0000;
      p30_uge_6683 <= 1'h0;
      p30_bivisor__1 <= 33'h0_0000_0000;
      p30_uge_6691 <= 1'h0;
      p30_uge_6771 <= 1'h0;
      p30_uge_6851 <= 1'h0;
      p30_uge_6931 <= 1'h0;
      p30_uge_7011 <= 1'h0;
      p30_uge_7091 <= 1'h0;
      p30_uge_7171 <= 1'h0;
      p30_uge_7251 <= 1'h0;
      p30_uge_7331 <= 1'h0;
      p30_uge_7411 <= 1'h0;
      p30_uge_7491 <= 1'h0;
      p30_uge_7571 <= 1'h0;
      p30_uge_7651 <= 1'h0;
      p30_uge_7731 <= 1'h0;
      p30_uge_7811 <= 1'h0;
      p30_uge_7891 <= 1'h0;
      p30_uge_7971 <= 1'h0;
      p30_uge_8051 <= 1'h0;
      p30_uge_8131 <= 1'h0;
      p30_uge_8211 <= 1'h0;
      p30_uge_8291 <= 1'h0;
      p30_uge_8371 <= 1'h0;
      p30_uge_8451 <= 1'h0;
      p30_uge_8531 <= 1'h0;
      p30_uge_8611 <= 1'h0;
      p30_uge_8691 <= 1'h0;
      p30_uge_8771 <= 1'h0;
      p30_uge_8851 <= 1'h0;
      p30_uge_8931 <= 1'h0;
      p30_concat_9010 <= 32'h0000_0000;
      p30_uge_9011 <= 1'h0;
      p30_bit_slice_6607 <= 1'h0;
      p30_negated <= 1'h0;
      p31_uge_6683 <= 1'h0;
      p31_uge_6691 <= 1'h0;
      p31_uge_6771 <= 1'h0;
      p31_uge_6851 <= 1'h0;
      p31_uge_6931 <= 1'h0;
      p31_uge_7011 <= 1'h0;
      p31_uge_7091 <= 1'h0;
      p31_uge_7171 <= 1'h0;
      p31_uge_7251 <= 1'h0;
      p31_uge_7331 <= 1'h0;
      p31_uge_7411 <= 1'h0;
      p31_uge_7491 <= 1'h0;
      p31_uge_7571 <= 1'h0;
      p31_uge_7651 <= 1'h0;
      p31_uge_7731 <= 1'h0;
      p31_uge_7811 <= 1'h0;
      p31_uge_7891 <= 1'h0;
      p31_uge_7971 <= 1'h0;
      p31_uge_8051 <= 1'h0;
      p31_uge_8131 <= 1'h0;
      p31_uge_8211 <= 1'h0;
      p31_uge_8291 <= 1'h0;
      p31_uge_8371 <= 1'h0;
      p31_uge_8451 <= 1'h0;
      p31_uge_8531 <= 1'h0;
      p31_uge_8611 <= 1'h0;
      p31_uge_8691 <= 1'h0;
      p31_uge_8771 <= 1'h0;
      p31_uge_8851 <= 1'h0;
      p31_uge_8931 <= 1'h0;
      p31_uge_9011 <= 1'h0;
      p31_q__32_squeezed_portion_0_width_1 <= 1'h0;
      p31_negated <= 1'h0;
      p0_valid <= 1'h0;
      p1_valid <= 1'h0;
      p2_valid <= 1'h0;
      p3_valid <= 1'h0;
      p4_valid <= 1'h0;
      p5_valid <= 1'h0;
      p6_valid <= 1'h0;
      p7_valid <= 1'h0;
      p8_valid <= 1'h0;
      p9_valid <= 1'h0;
      p10_valid <= 1'h0;
      p11_valid <= 1'h0;
      p12_valid <= 1'h0;
      p13_valid <= 1'h0;
      p14_valid <= 1'h0;
      p15_valid <= 1'h0;
      p16_valid <= 1'h0;
      p17_valid <= 1'h0;
      p18_valid <= 1'h0;
      p19_valid <= 1'h0;
      p20_valid <= 1'h0;
      p21_valid <= 1'h0;
      p22_valid <= 1'h0;
      p23_valid <= 1'h0;
      p24_valid <= 1'h0;
      p25_valid <= 1'h0;
      p26_valid <= 1'h0;
      p27_valid <= 1'h0;
      p28_valid <= 1'h0;
      p29_valid <= 1'h0;
      p30_valid <= 1'h0;
      p31_valid <= 1'h0;
      p32_valid <= 1'h0;
      p33_valid <= 1'h0;
      p34_valid <= 1'h0;
      __xls_float_ips__result_reg <= 32'h0000_0000;
      __xls_float_ips__result_valid_reg <= 1'h0;
    end else begin
      p0_concat_6575 <= p0_data_enable ? concat_6575 : p0_concat_6575;
      p0_b <= p0_data_enable ? xls_float_ips__rhs : p0_b;
      p0_bit_slice_6577 <= p0_data_enable ? bit_slice_6577 : p0_bit_slice_6577;
      p0_bit_slice_6578 <= p0_data_enable ? bit_slice_6578 : p0_bit_slice_6578;
      p0_bit_slice_6579 <= p0_data_enable ? bit_slice_6579 : p0_bit_slice_6579;
      p0_bit_slice_6580 <= p0_data_enable ? bit_slice_6580 : p0_bit_slice_6580;
      p0_bit_slice_6581 <= p0_data_enable ? bit_slice_6581 : p0_bit_slice_6581;
      p0_bit_slice_6582 <= p0_data_enable ? bit_slice_6582 : p0_bit_slice_6582;
      p0_bit_slice_6583 <= p0_data_enable ? bit_slice_6583 : p0_bit_slice_6583;
      p0_bit_slice_6584 <= p0_data_enable ? bit_slice_6584 : p0_bit_slice_6584;
      p0_bit_slice_6585 <= p0_data_enable ? bit_slice_6585 : p0_bit_slice_6585;
      p0_bit_slice_6586 <= p0_data_enable ? bit_slice_6586 : p0_bit_slice_6586;
      p0_bit_slice_6587 <= p0_data_enable ? bit_slice_6587 : p0_bit_slice_6587;
      p0_bit_slice_6588 <= p0_data_enable ? bit_slice_6588 : p0_bit_slice_6588;
      p0_bit_slice_6589 <= p0_data_enable ? bit_slice_6589 : p0_bit_slice_6589;
      p0_bit_slice_6590 <= p0_data_enable ? bit_slice_6590 : p0_bit_slice_6590;
      p0_bit_slice_6591 <= p0_data_enable ? bit_slice_6591 : p0_bit_slice_6591;
      p0_bit_slice_6592 <= p0_data_enable ? bit_slice_6592 : p0_bit_slice_6592;
      p0_bit_slice_6593 <= p0_data_enable ? bit_slice_6593 : p0_bit_slice_6593;
      p0_bit_slice_6594 <= p0_data_enable ? bit_slice_6594 : p0_bit_slice_6594;
      p0_bit_slice_6595 <= p0_data_enable ? bit_slice_6595 : p0_bit_slice_6595;
      p0_bit_slice_6596 <= p0_data_enable ? bit_slice_6596 : p0_bit_slice_6596;
      p0_bit_slice_6597 <= p0_data_enable ? bit_slice_6597 : p0_bit_slice_6597;
      p0_bit_slice_6598 <= p0_data_enable ? bit_slice_6598 : p0_bit_slice_6598;
      p0_bit_slice_6599 <= p0_data_enable ? bit_slice_6599 : p0_bit_slice_6599;
      p0_bit_slice_6600 <= p0_data_enable ? bit_slice_6600 : p0_bit_slice_6600;
      p0_bit_slice_6601 <= p0_data_enable ? bit_slice_6601 : p0_bit_slice_6601;
      p0_bit_slice_6602 <= p0_data_enable ? bit_slice_6602 : p0_bit_slice_6602;
      p0_bit_slice_6603 <= p0_data_enable ? bit_slice_6603 : p0_bit_slice_6603;
      p0_bit_slice_6604 <= p0_data_enable ? bit_slice_6604 : p0_bit_slice_6604;
      p0_bit_slice_6605 <= p0_data_enable ? bit_slice_6605 : p0_bit_slice_6605;
      p0_bit_slice_6606 <= p0_data_enable ? bit_slice_6606 : p0_bit_slice_6606;
      p0_bit_slice_6607 <= p0_data_enable ? bit_slice_6607 : p0_bit_slice_6607;
      p0_negated <= p0_data_enable ? negated : p0_negated;
      p1_b <= p1_data_enable ? p0_b : p1_b;
      p1_uge_6683 <= p1_data_enable ? uge_6683 : p1_uge_6683;
      p1_bivisor__1 <= p1_data_enable ? bivisor__1 : p1_bivisor__1;
      p1_concat_6690 <= p1_data_enable ? concat_6690 : p1_concat_6690;
      p1_uge_6691 <= p1_data_enable ? uge_6691 : p1_uge_6691;
      p1_bit_slice_6578 <= p1_data_enable ? p0_bit_slice_6578 : p1_bit_slice_6578;
      p1_bit_slice_6579 <= p1_data_enable ? p0_bit_slice_6579 : p1_bit_slice_6579;
      p1_bit_slice_6580 <= p1_data_enable ? p0_bit_slice_6580 : p1_bit_slice_6580;
      p1_bit_slice_6581 <= p1_data_enable ? p0_bit_slice_6581 : p1_bit_slice_6581;
      p1_bit_slice_6582 <= p1_data_enable ? p0_bit_slice_6582 : p1_bit_slice_6582;
      p1_bit_slice_6583 <= p1_data_enable ? p0_bit_slice_6583 : p1_bit_slice_6583;
      p1_bit_slice_6584 <= p1_data_enable ? p0_bit_slice_6584 : p1_bit_slice_6584;
      p1_bit_slice_6585 <= p1_data_enable ? p0_bit_slice_6585 : p1_bit_slice_6585;
      p1_bit_slice_6586 <= p1_data_enable ? p0_bit_slice_6586 : p1_bit_slice_6586;
      p1_bit_slice_6587 <= p1_data_enable ? p0_bit_slice_6587 : p1_bit_slice_6587;
      p1_bit_slice_6588 <= p1_data_enable ? p0_bit_slice_6588 : p1_bit_slice_6588;
      p1_bit_slice_6589 <= p1_data_enable ? p0_bit_slice_6589 : p1_bit_slice_6589;
      p1_bit_slice_6590 <= p1_data_enable ? p0_bit_slice_6590 : p1_bit_slice_6590;
      p1_bit_slice_6591 <= p1_data_enable ? p0_bit_slice_6591 : p1_bit_slice_6591;
      p1_bit_slice_6592 <= p1_data_enable ? p0_bit_slice_6592 : p1_bit_slice_6592;
      p1_bit_slice_6593 <= p1_data_enable ? p0_bit_slice_6593 : p1_bit_slice_6593;
      p1_bit_slice_6594 <= p1_data_enable ? p0_bit_slice_6594 : p1_bit_slice_6594;
      p1_bit_slice_6595 <= p1_data_enable ? p0_bit_slice_6595 : p1_bit_slice_6595;
      p1_bit_slice_6596 <= p1_data_enable ? p0_bit_slice_6596 : p1_bit_slice_6596;
      p1_bit_slice_6597 <= p1_data_enable ? p0_bit_slice_6597 : p1_bit_slice_6597;
      p1_bit_slice_6598 <= p1_data_enable ? p0_bit_slice_6598 : p1_bit_slice_6598;
      p1_bit_slice_6599 <= p1_data_enable ? p0_bit_slice_6599 : p1_bit_slice_6599;
      p1_bit_slice_6600 <= p1_data_enable ? p0_bit_slice_6600 : p1_bit_slice_6600;
      p1_bit_slice_6601 <= p1_data_enable ? p0_bit_slice_6601 : p1_bit_slice_6601;
      p1_bit_slice_6602 <= p1_data_enable ? p0_bit_slice_6602 : p1_bit_slice_6602;
      p1_bit_slice_6603 <= p1_data_enable ? p0_bit_slice_6603 : p1_bit_slice_6603;
      p1_bit_slice_6604 <= p1_data_enable ? p0_bit_slice_6604 : p1_bit_slice_6604;
      p1_bit_slice_6605 <= p1_data_enable ? p0_bit_slice_6605 : p1_bit_slice_6605;
      p1_bit_slice_6606 <= p1_data_enable ? p0_bit_slice_6606 : p1_bit_slice_6606;
      p1_bit_slice_6607 <= p1_data_enable ? p0_bit_slice_6607 : p1_bit_slice_6607;
      p1_negated <= p1_data_enable ? p0_negated : p1_negated;
      p2_b <= p2_data_enable ? p1_b : p2_b;
      p2_uge_6683 <= p2_data_enable ? p1_uge_6683 : p2_uge_6683;
      p2_bivisor__1 <= p2_data_enable ? p1_bivisor__1 : p2_bivisor__1;
      p2_uge_6691 <= p2_data_enable ? p1_uge_6691 : p2_uge_6691;
      p2_concat_6770 <= p2_data_enable ? concat_6770 : p2_concat_6770;
      p2_uge_6771 <= p2_data_enable ? uge_6771 : p2_uge_6771;
      p2_bit_slice_6579 <= p2_data_enable ? p1_bit_slice_6579 : p2_bit_slice_6579;
      p2_bit_slice_6580 <= p2_data_enable ? p1_bit_slice_6580 : p2_bit_slice_6580;
      p2_bit_slice_6581 <= p2_data_enable ? p1_bit_slice_6581 : p2_bit_slice_6581;
      p2_bit_slice_6582 <= p2_data_enable ? p1_bit_slice_6582 : p2_bit_slice_6582;
      p2_bit_slice_6583 <= p2_data_enable ? p1_bit_slice_6583 : p2_bit_slice_6583;
      p2_bit_slice_6584 <= p2_data_enable ? p1_bit_slice_6584 : p2_bit_slice_6584;
      p2_bit_slice_6585 <= p2_data_enable ? p1_bit_slice_6585 : p2_bit_slice_6585;
      p2_bit_slice_6586 <= p2_data_enable ? p1_bit_slice_6586 : p2_bit_slice_6586;
      p2_bit_slice_6587 <= p2_data_enable ? p1_bit_slice_6587 : p2_bit_slice_6587;
      p2_bit_slice_6588 <= p2_data_enable ? p1_bit_slice_6588 : p2_bit_slice_6588;
      p2_bit_slice_6589 <= p2_data_enable ? p1_bit_slice_6589 : p2_bit_slice_6589;
      p2_bit_slice_6590 <= p2_data_enable ? p1_bit_slice_6590 : p2_bit_slice_6590;
      p2_bit_slice_6591 <= p2_data_enable ? p1_bit_slice_6591 : p2_bit_slice_6591;
      p2_bit_slice_6592 <= p2_data_enable ? p1_bit_slice_6592 : p2_bit_slice_6592;
      p2_bit_slice_6593 <= p2_data_enable ? p1_bit_slice_6593 : p2_bit_slice_6593;
      p2_bit_slice_6594 <= p2_data_enable ? p1_bit_slice_6594 : p2_bit_slice_6594;
      p2_bit_slice_6595 <= p2_data_enable ? p1_bit_slice_6595 : p2_bit_slice_6595;
      p2_bit_slice_6596 <= p2_data_enable ? p1_bit_slice_6596 : p2_bit_slice_6596;
      p2_bit_slice_6597 <= p2_data_enable ? p1_bit_slice_6597 : p2_bit_slice_6597;
      p2_bit_slice_6598 <= p2_data_enable ? p1_bit_slice_6598 : p2_bit_slice_6598;
      p2_bit_slice_6599 <= p2_data_enable ? p1_bit_slice_6599 : p2_bit_slice_6599;
      p2_bit_slice_6600 <= p2_data_enable ? p1_bit_slice_6600 : p2_bit_slice_6600;
      p2_bit_slice_6601 <= p2_data_enable ? p1_bit_slice_6601 : p2_bit_slice_6601;
      p2_bit_slice_6602 <= p2_data_enable ? p1_bit_slice_6602 : p2_bit_slice_6602;
      p2_bit_slice_6603 <= p2_data_enable ? p1_bit_slice_6603 : p2_bit_slice_6603;
      p2_bit_slice_6604 <= p2_data_enable ? p1_bit_slice_6604 : p2_bit_slice_6604;
      p2_bit_slice_6605 <= p2_data_enable ? p1_bit_slice_6605 : p2_bit_slice_6605;
      p2_bit_slice_6606 <= p2_data_enable ? p1_bit_slice_6606 : p2_bit_slice_6606;
      p2_bit_slice_6607 <= p2_data_enable ? p1_bit_slice_6607 : p2_bit_slice_6607;
      p2_negated <= p2_data_enable ? p1_negated : p2_negated;
      p3_b <= p3_data_enable ? p2_b : p3_b;
      p3_uge_6683 <= p3_data_enable ? p2_uge_6683 : p3_uge_6683;
      p3_bivisor__1 <= p3_data_enable ? p2_bivisor__1 : p3_bivisor__1;
      p3_uge_6691 <= p3_data_enable ? p2_uge_6691 : p3_uge_6691;
      p3_uge_6771 <= p3_data_enable ? p2_uge_6771 : p3_uge_6771;
      p3_concat_6850 <= p3_data_enable ? concat_6850 : p3_concat_6850;
      p3_uge_6851 <= p3_data_enable ? uge_6851 : p3_uge_6851;
      p3_bit_slice_6580 <= p3_data_enable ? p2_bit_slice_6580 : p3_bit_slice_6580;
      p3_bit_slice_6581 <= p3_data_enable ? p2_bit_slice_6581 : p3_bit_slice_6581;
      p3_bit_slice_6582 <= p3_data_enable ? p2_bit_slice_6582 : p3_bit_slice_6582;
      p3_bit_slice_6583 <= p3_data_enable ? p2_bit_slice_6583 : p3_bit_slice_6583;
      p3_bit_slice_6584 <= p3_data_enable ? p2_bit_slice_6584 : p3_bit_slice_6584;
      p3_bit_slice_6585 <= p3_data_enable ? p2_bit_slice_6585 : p3_bit_slice_6585;
      p3_bit_slice_6586 <= p3_data_enable ? p2_bit_slice_6586 : p3_bit_slice_6586;
      p3_bit_slice_6587 <= p3_data_enable ? p2_bit_slice_6587 : p3_bit_slice_6587;
      p3_bit_slice_6588 <= p3_data_enable ? p2_bit_slice_6588 : p3_bit_slice_6588;
      p3_bit_slice_6589 <= p3_data_enable ? p2_bit_slice_6589 : p3_bit_slice_6589;
      p3_bit_slice_6590 <= p3_data_enable ? p2_bit_slice_6590 : p3_bit_slice_6590;
      p3_bit_slice_6591 <= p3_data_enable ? p2_bit_slice_6591 : p3_bit_slice_6591;
      p3_bit_slice_6592 <= p3_data_enable ? p2_bit_slice_6592 : p3_bit_slice_6592;
      p3_bit_slice_6593 <= p3_data_enable ? p2_bit_slice_6593 : p3_bit_slice_6593;
      p3_bit_slice_6594 <= p3_data_enable ? p2_bit_slice_6594 : p3_bit_slice_6594;
      p3_bit_slice_6595 <= p3_data_enable ? p2_bit_slice_6595 : p3_bit_slice_6595;
      p3_bit_slice_6596 <= p3_data_enable ? p2_bit_slice_6596 : p3_bit_slice_6596;
      p3_bit_slice_6597 <= p3_data_enable ? p2_bit_slice_6597 : p3_bit_slice_6597;
      p3_bit_slice_6598 <= p3_data_enable ? p2_bit_slice_6598 : p3_bit_slice_6598;
      p3_bit_slice_6599 <= p3_data_enable ? p2_bit_slice_6599 : p3_bit_slice_6599;
      p3_bit_slice_6600 <= p3_data_enable ? p2_bit_slice_6600 : p3_bit_slice_6600;
      p3_bit_slice_6601 <= p3_data_enable ? p2_bit_slice_6601 : p3_bit_slice_6601;
      p3_bit_slice_6602 <= p3_data_enable ? p2_bit_slice_6602 : p3_bit_slice_6602;
      p3_bit_slice_6603 <= p3_data_enable ? p2_bit_slice_6603 : p3_bit_slice_6603;
      p3_bit_slice_6604 <= p3_data_enable ? p2_bit_slice_6604 : p3_bit_slice_6604;
      p3_bit_slice_6605 <= p3_data_enable ? p2_bit_slice_6605 : p3_bit_slice_6605;
      p3_bit_slice_6606 <= p3_data_enable ? p2_bit_slice_6606 : p3_bit_slice_6606;
      p3_bit_slice_6607 <= p3_data_enable ? p2_bit_slice_6607 : p3_bit_slice_6607;
      p3_negated <= p3_data_enable ? p2_negated : p3_negated;
      p4_b <= p4_data_enable ? p3_b : p4_b;
      p4_uge_6683 <= p4_data_enable ? p3_uge_6683 : p4_uge_6683;
      p4_bivisor__1 <= p4_data_enable ? p3_bivisor__1 : p4_bivisor__1;
      p4_uge_6691 <= p4_data_enable ? p3_uge_6691 : p4_uge_6691;
      p4_uge_6771 <= p4_data_enable ? p3_uge_6771 : p4_uge_6771;
      p4_uge_6851 <= p4_data_enable ? p3_uge_6851 : p4_uge_6851;
      p4_concat_6930 <= p4_data_enable ? concat_6930 : p4_concat_6930;
      p4_uge_6931 <= p4_data_enable ? uge_6931 : p4_uge_6931;
      p4_bit_slice_6581 <= p4_data_enable ? p3_bit_slice_6581 : p4_bit_slice_6581;
      p4_bit_slice_6582 <= p4_data_enable ? p3_bit_slice_6582 : p4_bit_slice_6582;
      p4_bit_slice_6583 <= p4_data_enable ? p3_bit_slice_6583 : p4_bit_slice_6583;
      p4_bit_slice_6584 <= p4_data_enable ? p3_bit_slice_6584 : p4_bit_slice_6584;
      p4_bit_slice_6585 <= p4_data_enable ? p3_bit_slice_6585 : p4_bit_slice_6585;
      p4_bit_slice_6586 <= p4_data_enable ? p3_bit_slice_6586 : p4_bit_slice_6586;
      p4_bit_slice_6587 <= p4_data_enable ? p3_bit_slice_6587 : p4_bit_slice_6587;
      p4_bit_slice_6588 <= p4_data_enable ? p3_bit_slice_6588 : p4_bit_slice_6588;
      p4_bit_slice_6589 <= p4_data_enable ? p3_bit_slice_6589 : p4_bit_slice_6589;
      p4_bit_slice_6590 <= p4_data_enable ? p3_bit_slice_6590 : p4_bit_slice_6590;
      p4_bit_slice_6591 <= p4_data_enable ? p3_bit_slice_6591 : p4_bit_slice_6591;
      p4_bit_slice_6592 <= p4_data_enable ? p3_bit_slice_6592 : p4_bit_slice_6592;
      p4_bit_slice_6593 <= p4_data_enable ? p3_bit_slice_6593 : p4_bit_slice_6593;
      p4_bit_slice_6594 <= p4_data_enable ? p3_bit_slice_6594 : p4_bit_slice_6594;
      p4_bit_slice_6595 <= p4_data_enable ? p3_bit_slice_6595 : p4_bit_slice_6595;
      p4_bit_slice_6596 <= p4_data_enable ? p3_bit_slice_6596 : p4_bit_slice_6596;
      p4_bit_slice_6597 <= p4_data_enable ? p3_bit_slice_6597 : p4_bit_slice_6597;
      p4_bit_slice_6598 <= p4_data_enable ? p3_bit_slice_6598 : p4_bit_slice_6598;
      p4_bit_slice_6599 <= p4_data_enable ? p3_bit_slice_6599 : p4_bit_slice_6599;
      p4_bit_slice_6600 <= p4_data_enable ? p3_bit_slice_6600 : p4_bit_slice_6600;
      p4_bit_slice_6601 <= p4_data_enable ? p3_bit_slice_6601 : p4_bit_slice_6601;
      p4_bit_slice_6602 <= p4_data_enable ? p3_bit_slice_6602 : p4_bit_slice_6602;
      p4_bit_slice_6603 <= p4_data_enable ? p3_bit_slice_6603 : p4_bit_slice_6603;
      p4_bit_slice_6604 <= p4_data_enable ? p3_bit_slice_6604 : p4_bit_slice_6604;
      p4_bit_slice_6605 <= p4_data_enable ? p3_bit_slice_6605 : p4_bit_slice_6605;
      p4_bit_slice_6606 <= p4_data_enable ? p3_bit_slice_6606 : p4_bit_slice_6606;
      p4_bit_slice_6607 <= p4_data_enable ? p3_bit_slice_6607 : p4_bit_slice_6607;
      p4_negated <= p4_data_enable ? p3_negated : p4_negated;
      p5_b <= p5_data_enable ? p4_b : p5_b;
      p5_uge_6683 <= p5_data_enable ? p4_uge_6683 : p5_uge_6683;
      p5_bivisor__1 <= p5_data_enable ? p4_bivisor__1 : p5_bivisor__1;
      p5_uge_6691 <= p5_data_enable ? p4_uge_6691 : p5_uge_6691;
      p5_uge_6771 <= p5_data_enable ? p4_uge_6771 : p5_uge_6771;
      p5_uge_6851 <= p5_data_enable ? p4_uge_6851 : p5_uge_6851;
      p5_uge_6931 <= p5_data_enable ? p4_uge_6931 : p5_uge_6931;
      p5_concat_7010 <= p5_data_enable ? concat_7010 : p5_concat_7010;
      p5_uge_7011 <= p5_data_enable ? uge_7011 : p5_uge_7011;
      p5_bit_slice_6582 <= p5_data_enable ? p4_bit_slice_6582 : p5_bit_slice_6582;
      p5_bit_slice_6583 <= p5_data_enable ? p4_bit_slice_6583 : p5_bit_slice_6583;
      p5_bit_slice_6584 <= p5_data_enable ? p4_bit_slice_6584 : p5_bit_slice_6584;
      p5_bit_slice_6585 <= p5_data_enable ? p4_bit_slice_6585 : p5_bit_slice_6585;
      p5_bit_slice_6586 <= p5_data_enable ? p4_bit_slice_6586 : p5_bit_slice_6586;
      p5_bit_slice_6587 <= p5_data_enable ? p4_bit_slice_6587 : p5_bit_slice_6587;
      p5_bit_slice_6588 <= p5_data_enable ? p4_bit_slice_6588 : p5_bit_slice_6588;
      p5_bit_slice_6589 <= p5_data_enable ? p4_bit_slice_6589 : p5_bit_slice_6589;
      p5_bit_slice_6590 <= p5_data_enable ? p4_bit_slice_6590 : p5_bit_slice_6590;
      p5_bit_slice_6591 <= p5_data_enable ? p4_bit_slice_6591 : p5_bit_slice_6591;
      p5_bit_slice_6592 <= p5_data_enable ? p4_bit_slice_6592 : p5_bit_slice_6592;
      p5_bit_slice_6593 <= p5_data_enable ? p4_bit_slice_6593 : p5_bit_slice_6593;
      p5_bit_slice_6594 <= p5_data_enable ? p4_bit_slice_6594 : p5_bit_slice_6594;
      p5_bit_slice_6595 <= p5_data_enable ? p4_bit_slice_6595 : p5_bit_slice_6595;
      p5_bit_slice_6596 <= p5_data_enable ? p4_bit_slice_6596 : p5_bit_slice_6596;
      p5_bit_slice_6597 <= p5_data_enable ? p4_bit_slice_6597 : p5_bit_slice_6597;
      p5_bit_slice_6598 <= p5_data_enable ? p4_bit_slice_6598 : p5_bit_slice_6598;
      p5_bit_slice_6599 <= p5_data_enable ? p4_bit_slice_6599 : p5_bit_slice_6599;
      p5_bit_slice_6600 <= p5_data_enable ? p4_bit_slice_6600 : p5_bit_slice_6600;
      p5_bit_slice_6601 <= p5_data_enable ? p4_bit_slice_6601 : p5_bit_slice_6601;
      p5_bit_slice_6602 <= p5_data_enable ? p4_bit_slice_6602 : p5_bit_slice_6602;
      p5_bit_slice_6603 <= p5_data_enable ? p4_bit_slice_6603 : p5_bit_slice_6603;
      p5_bit_slice_6604 <= p5_data_enable ? p4_bit_slice_6604 : p5_bit_slice_6604;
      p5_bit_slice_6605 <= p5_data_enable ? p4_bit_slice_6605 : p5_bit_slice_6605;
      p5_bit_slice_6606 <= p5_data_enable ? p4_bit_slice_6606 : p5_bit_slice_6606;
      p5_bit_slice_6607 <= p5_data_enable ? p4_bit_slice_6607 : p5_bit_slice_6607;
      p5_negated <= p5_data_enable ? p4_negated : p5_negated;
      p6_b <= p6_data_enable ? p5_b : p6_b;
      p6_uge_6683 <= p6_data_enable ? p5_uge_6683 : p6_uge_6683;
      p6_bivisor__1 <= p6_data_enable ? p5_bivisor__1 : p6_bivisor__1;
      p6_uge_6691 <= p6_data_enable ? p5_uge_6691 : p6_uge_6691;
      p6_uge_6771 <= p6_data_enable ? p5_uge_6771 : p6_uge_6771;
      p6_uge_6851 <= p6_data_enable ? p5_uge_6851 : p6_uge_6851;
      p6_uge_6931 <= p6_data_enable ? p5_uge_6931 : p6_uge_6931;
      p6_uge_7011 <= p6_data_enable ? p5_uge_7011 : p6_uge_7011;
      p6_concat_7090 <= p6_data_enable ? concat_7090 : p6_concat_7090;
      p6_uge_7091 <= p6_data_enable ? uge_7091 : p6_uge_7091;
      p6_bit_slice_6583 <= p6_data_enable ? p5_bit_slice_6583 : p6_bit_slice_6583;
      p6_bit_slice_6584 <= p6_data_enable ? p5_bit_slice_6584 : p6_bit_slice_6584;
      p6_bit_slice_6585 <= p6_data_enable ? p5_bit_slice_6585 : p6_bit_slice_6585;
      p6_bit_slice_6586 <= p6_data_enable ? p5_bit_slice_6586 : p6_bit_slice_6586;
      p6_bit_slice_6587 <= p6_data_enable ? p5_bit_slice_6587 : p6_bit_slice_6587;
      p6_bit_slice_6588 <= p6_data_enable ? p5_bit_slice_6588 : p6_bit_slice_6588;
      p6_bit_slice_6589 <= p6_data_enable ? p5_bit_slice_6589 : p6_bit_slice_6589;
      p6_bit_slice_6590 <= p6_data_enable ? p5_bit_slice_6590 : p6_bit_slice_6590;
      p6_bit_slice_6591 <= p6_data_enable ? p5_bit_slice_6591 : p6_bit_slice_6591;
      p6_bit_slice_6592 <= p6_data_enable ? p5_bit_slice_6592 : p6_bit_slice_6592;
      p6_bit_slice_6593 <= p6_data_enable ? p5_bit_slice_6593 : p6_bit_slice_6593;
      p6_bit_slice_6594 <= p6_data_enable ? p5_bit_slice_6594 : p6_bit_slice_6594;
      p6_bit_slice_6595 <= p6_data_enable ? p5_bit_slice_6595 : p6_bit_slice_6595;
      p6_bit_slice_6596 <= p6_data_enable ? p5_bit_slice_6596 : p6_bit_slice_6596;
      p6_bit_slice_6597 <= p6_data_enable ? p5_bit_slice_6597 : p6_bit_slice_6597;
      p6_bit_slice_6598 <= p6_data_enable ? p5_bit_slice_6598 : p6_bit_slice_6598;
      p6_bit_slice_6599 <= p6_data_enable ? p5_bit_slice_6599 : p6_bit_slice_6599;
      p6_bit_slice_6600 <= p6_data_enable ? p5_bit_slice_6600 : p6_bit_slice_6600;
      p6_bit_slice_6601 <= p6_data_enable ? p5_bit_slice_6601 : p6_bit_slice_6601;
      p6_bit_slice_6602 <= p6_data_enable ? p5_bit_slice_6602 : p6_bit_slice_6602;
      p6_bit_slice_6603 <= p6_data_enable ? p5_bit_slice_6603 : p6_bit_slice_6603;
      p6_bit_slice_6604 <= p6_data_enable ? p5_bit_slice_6604 : p6_bit_slice_6604;
      p6_bit_slice_6605 <= p6_data_enable ? p5_bit_slice_6605 : p6_bit_slice_6605;
      p6_bit_slice_6606 <= p6_data_enable ? p5_bit_slice_6606 : p6_bit_slice_6606;
      p6_bit_slice_6607 <= p6_data_enable ? p5_bit_slice_6607 : p6_bit_slice_6607;
      p6_negated <= p6_data_enable ? p5_negated : p6_negated;
      p7_b <= p7_data_enable ? p6_b : p7_b;
      p7_uge_6683 <= p7_data_enable ? p6_uge_6683 : p7_uge_6683;
      p7_bivisor__1 <= p7_data_enable ? p6_bivisor__1 : p7_bivisor__1;
      p7_uge_6691 <= p7_data_enable ? p6_uge_6691 : p7_uge_6691;
      p7_uge_6771 <= p7_data_enable ? p6_uge_6771 : p7_uge_6771;
      p7_uge_6851 <= p7_data_enable ? p6_uge_6851 : p7_uge_6851;
      p7_uge_6931 <= p7_data_enable ? p6_uge_6931 : p7_uge_6931;
      p7_uge_7011 <= p7_data_enable ? p6_uge_7011 : p7_uge_7011;
      p7_uge_7091 <= p7_data_enable ? p6_uge_7091 : p7_uge_7091;
      p7_concat_7170 <= p7_data_enable ? concat_7170 : p7_concat_7170;
      p7_uge_7171 <= p7_data_enable ? uge_7171 : p7_uge_7171;
      p7_bit_slice_6584 <= p7_data_enable ? p6_bit_slice_6584 : p7_bit_slice_6584;
      p7_bit_slice_6585 <= p7_data_enable ? p6_bit_slice_6585 : p7_bit_slice_6585;
      p7_bit_slice_6586 <= p7_data_enable ? p6_bit_slice_6586 : p7_bit_slice_6586;
      p7_bit_slice_6587 <= p7_data_enable ? p6_bit_slice_6587 : p7_bit_slice_6587;
      p7_bit_slice_6588 <= p7_data_enable ? p6_bit_slice_6588 : p7_bit_slice_6588;
      p7_bit_slice_6589 <= p7_data_enable ? p6_bit_slice_6589 : p7_bit_slice_6589;
      p7_bit_slice_6590 <= p7_data_enable ? p6_bit_slice_6590 : p7_bit_slice_6590;
      p7_bit_slice_6591 <= p7_data_enable ? p6_bit_slice_6591 : p7_bit_slice_6591;
      p7_bit_slice_6592 <= p7_data_enable ? p6_bit_slice_6592 : p7_bit_slice_6592;
      p7_bit_slice_6593 <= p7_data_enable ? p6_bit_slice_6593 : p7_bit_slice_6593;
      p7_bit_slice_6594 <= p7_data_enable ? p6_bit_slice_6594 : p7_bit_slice_6594;
      p7_bit_slice_6595 <= p7_data_enable ? p6_bit_slice_6595 : p7_bit_slice_6595;
      p7_bit_slice_6596 <= p7_data_enable ? p6_bit_slice_6596 : p7_bit_slice_6596;
      p7_bit_slice_6597 <= p7_data_enable ? p6_bit_slice_6597 : p7_bit_slice_6597;
      p7_bit_slice_6598 <= p7_data_enable ? p6_bit_slice_6598 : p7_bit_slice_6598;
      p7_bit_slice_6599 <= p7_data_enable ? p6_bit_slice_6599 : p7_bit_slice_6599;
      p7_bit_slice_6600 <= p7_data_enable ? p6_bit_slice_6600 : p7_bit_slice_6600;
      p7_bit_slice_6601 <= p7_data_enable ? p6_bit_slice_6601 : p7_bit_slice_6601;
      p7_bit_slice_6602 <= p7_data_enable ? p6_bit_slice_6602 : p7_bit_slice_6602;
      p7_bit_slice_6603 <= p7_data_enable ? p6_bit_slice_6603 : p7_bit_slice_6603;
      p7_bit_slice_6604 <= p7_data_enable ? p6_bit_slice_6604 : p7_bit_slice_6604;
      p7_bit_slice_6605 <= p7_data_enable ? p6_bit_slice_6605 : p7_bit_slice_6605;
      p7_bit_slice_6606 <= p7_data_enable ? p6_bit_slice_6606 : p7_bit_slice_6606;
      p7_bit_slice_6607 <= p7_data_enable ? p6_bit_slice_6607 : p7_bit_slice_6607;
      p7_negated <= p7_data_enable ? p6_negated : p7_negated;
      p8_b <= p8_data_enable ? p7_b : p8_b;
      p8_uge_6683 <= p8_data_enable ? p7_uge_6683 : p8_uge_6683;
      p8_bivisor__1 <= p8_data_enable ? p7_bivisor__1 : p8_bivisor__1;
      p8_uge_6691 <= p8_data_enable ? p7_uge_6691 : p8_uge_6691;
      p8_uge_6771 <= p8_data_enable ? p7_uge_6771 : p8_uge_6771;
      p8_uge_6851 <= p8_data_enable ? p7_uge_6851 : p8_uge_6851;
      p8_uge_6931 <= p8_data_enable ? p7_uge_6931 : p8_uge_6931;
      p8_uge_7011 <= p8_data_enable ? p7_uge_7011 : p8_uge_7011;
      p8_uge_7091 <= p8_data_enable ? p7_uge_7091 : p8_uge_7091;
      p8_uge_7171 <= p8_data_enable ? p7_uge_7171 : p8_uge_7171;
      p8_concat_7250 <= p8_data_enable ? concat_7250 : p8_concat_7250;
      p8_uge_7251 <= p8_data_enable ? uge_7251 : p8_uge_7251;
      p8_bit_slice_6585 <= p8_data_enable ? p7_bit_slice_6585 : p8_bit_slice_6585;
      p8_bit_slice_6586 <= p8_data_enable ? p7_bit_slice_6586 : p8_bit_slice_6586;
      p8_bit_slice_6587 <= p8_data_enable ? p7_bit_slice_6587 : p8_bit_slice_6587;
      p8_bit_slice_6588 <= p8_data_enable ? p7_bit_slice_6588 : p8_bit_slice_6588;
      p8_bit_slice_6589 <= p8_data_enable ? p7_bit_slice_6589 : p8_bit_slice_6589;
      p8_bit_slice_6590 <= p8_data_enable ? p7_bit_slice_6590 : p8_bit_slice_6590;
      p8_bit_slice_6591 <= p8_data_enable ? p7_bit_slice_6591 : p8_bit_slice_6591;
      p8_bit_slice_6592 <= p8_data_enable ? p7_bit_slice_6592 : p8_bit_slice_6592;
      p8_bit_slice_6593 <= p8_data_enable ? p7_bit_slice_6593 : p8_bit_slice_6593;
      p8_bit_slice_6594 <= p8_data_enable ? p7_bit_slice_6594 : p8_bit_slice_6594;
      p8_bit_slice_6595 <= p8_data_enable ? p7_bit_slice_6595 : p8_bit_slice_6595;
      p8_bit_slice_6596 <= p8_data_enable ? p7_bit_slice_6596 : p8_bit_slice_6596;
      p8_bit_slice_6597 <= p8_data_enable ? p7_bit_slice_6597 : p8_bit_slice_6597;
      p8_bit_slice_6598 <= p8_data_enable ? p7_bit_slice_6598 : p8_bit_slice_6598;
      p8_bit_slice_6599 <= p8_data_enable ? p7_bit_slice_6599 : p8_bit_slice_6599;
      p8_bit_slice_6600 <= p8_data_enable ? p7_bit_slice_6600 : p8_bit_slice_6600;
      p8_bit_slice_6601 <= p8_data_enable ? p7_bit_slice_6601 : p8_bit_slice_6601;
      p8_bit_slice_6602 <= p8_data_enable ? p7_bit_slice_6602 : p8_bit_slice_6602;
      p8_bit_slice_6603 <= p8_data_enable ? p7_bit_slice_6603 : p8_bit_slice_6603;
      p8_bit_slice_6604 <= p8_data_enable ? p7_bit_slice_6604 : p8_bit_slice_6604;
      p8_bit_slice_6605 <= p8_data_enable ? p7_bit_slice_6605 : p8_bit_slice_6605;
      p8_bit_slice_6606 <= p8_data_enable ? p7_bit_slice_6606 : p8_bit_slice_6606;
      p8_bit_slice_6607 <= p8_data_enable ? p7_bit_slice_6607 : p8_bit_slice_6607;
      p8_negated <= p8_data_enable ? p7_negated : p8_negated;
      p9_b <= p9_data_enable ? p8_b : p9_b;
      p9_uge_6683 <= p9_data_enable ? p8_uge_6683 : p9_uge_6683;
      p9_bivisor__1 <= p9_data_enable ? p8_bivisor__1 : p9_bivisor__1;
      p9_uge_6691 <= p9_data_enable ? p8_uge_6691 : p9_uge_6691;
      p9_uge_6771 <= p9_data_enable ? p8_uge_6771 : p9_uge_6771;
      p9_uge_6851 <= p9_data_enable ? p8_uge_6851 : p9_uge_6851;
      p9_uge_6931 <= p9_data_enable ? p8_uge_6931 : p9_uge_6931;
      p9_uge_7011 <= p9_data_enable ? p8_uge_7011 : p9_uge_7011;
      p9_uge_7091 <= p9_data_enable ? p8_uge_7091 : p9_uge_7091;
      p9_uge_7171 <= p9_data_enable ? p8_uge_7171 : p9_uge_7171;
      p9_uge_7251 <= p9_data_enable ? p8_uge_7251 : p9_uge_7251;
      p9_concat_7330 <= p9_data_enable ? concat_7330 : p9_concat_7330;
      p9_uge_7331 <= p9_data_enable ? uge_7331 : p9_uge_7331;
      p9_bit_slice_6586 <= p9_data_enable ? p8_bit_slice_6586 : p9_bit_slice_6586;
      p9_bit_slice_6587 <= p9_data_enable ? p8_bit_slice_6587 : p9_bit_slice_6587;
      p9_bit_slice_6588 <= p9_data_enable ? p8_bit_slice_6588 : p9_bit_slice_6588;
      p9_bit_slice_6589 <= p9_data_enable ? p8_bit_slice_6589 : p9_bit_slice_6589;
      p9_bit_slice_6590 <= p9_data_enable ? p8_bit_slice_6590 : p9_bit_slice_6590;
      p9_bit_slice_6591 <= p9_data_enable ? p8_bit_slice_6591 : p9_bit_slice_6591;
      p9_bit_slice_6592 <= p9_data_enable ? p8_bit_slice_6592 : p9_bit_slice_6592;
      p9_bit_slice_6593 <= p9_data_enable ? p8_bit_slice_6593 : p9_bit_slice_6593;
      p9_bit_slice_6594 <= p9_data_enable ? p8_bit_slice_6594 : p9_bit_slice_6594;
      p9_bit_slice_6595 <= p9_data_enable ? p8_bit_slice_6595 : p9_bit_slice_6595;
      p9_bit_slice_6596 <= p9_data_enable ? p8_bit_slice_6596 : p9_bit_slice_6596;
      p9_bit_slice_6597 <= p9_data_enable ? p8_bit_slice_6597 : p9_bit_slice_6597;
      p9_bit_slice_6598 <= p9_data_enable ? p8_bit_slice_6598 : p9_bit_slice_6598;
      p9_bit_slice_6599 <= p9_data_enable ? p8_bit_slice_6599 : p9_bit_slice_6599;
      p9_bit_slice_6600 <= p9_data_enable ? p8_bit_slice_6600 : p9_bit_slice_6600;
      p9_bit_slice_6601 <= p9_data_enable ? p8_bit_slice_6601 : p9_bit_slice_6601;
      p9_bit_slice_6602 <= p9_data_enable ? p8_bit_slice_6602 : p9_bit_slice_6602;
      p9_bit_slice_6603 <= p9_data_enable ? p8_bit_slice_6603 : p9_bit_slice_6603;
      p9_bit_slice_6604 <= p9_data_enable ? p8_bit_slice_6604 : p9_bit_slice_6604;
      p9_bit_slice_6605 <= p9_data_enable ? p8_bit_slice_6605 : p9_bit_slice_6605;
      p9_bit_slice_6606 <= p9_data_enable ? p8_bit_slice_6606 : p9_bit_slice_6606;
      p9_bit_slice_6607 <= p9_data_enable ? p8_bit_slice_6607 : p9_bit_slice_6607;
      p9_negated <= p9_data_enable ? p8_negated : p9_negated;
      p10_b <= p10_data_enable ? p9_b : p10_b;
      p10_uge_6683 <= p10_data_enable ? p9_uge_6683 : p10_uge_6683;
      p10_bivisor__1 <= p10_data_enable ? p9_bivisor__1 : p10_bivisor__1;
      p10_uge_6691 <= p10_data_enable ? p9_uge_6691 : p10_uge_6691;
      p10_uge_6771 <= p10_data_enable ? p9_uge_6771 : p10_uge_6771;
      p10_uge_6851 <= p10_data_enable ? p9_uge_6851 : p10_uge_6851;
      p10_uge_6931 <= p10_data_enable ? p9_uge_6931 : p10_uge_6931;
      p10_uge_7011 <= p10_data_enable ? p9_uge_7011 : p10_uge_7011;
      p10_uge_7091 <= p10_data_enable ? p9_uge_7091 : p10_uge_7091;
      p10_uge_7171 <= p10_data_enable ? p9_uge_7171 : p10_uge_7171;
      p10_uge_7251 <= p10_data_enable ? p9_uge_7251 : p10_uge_7251;
      p10_uge_7331 <= p10_data_enable ? p9_uge_7331 : p10_uge_7331;
      p10_concat_7410 <= p10_data_enable ? concat_7410 : p10_concat_7410;
      p10_uge_7411 <= p10_data_enable ? uge_7411 : p10_uge_7411;
      p10_bit_slice_6587 <= p10_data_enable ? p9_bit_slice_6587 : p10_bit_slice_6587;
      p10_bit_slice_6588 <= p10_data_enable ? p9_bit_slice_6588 : p10_bit_slice_6588;
      p10_bit_slice_6589 <= p10_data_enable ? p9_bit_slice_6589 : p10_bit_slice_6589;
      p10_bit_slice_6590 <= p10_data_enable ? p9_bit_slice_6590 : p10_bit_slice_6590;
      p10_bit_slice_6591 <= p10_data_enable ? p9_bit_slice_6591 : p10_bit_slice_6591;
      p10_bit_slice_6592 <= p10_data_enable ? p9_bit_slice_6592 : p10_bit_slice_6592;
      p10_bit_slice_6593 <= p10_data_enable ? p9_bit_slice_6593 : p10_bit_slice_6593;
      p10_bit_slice_6594 <= p10_data_enable ? p9_bit_slice_6594 : p10_bit_slice_6594;
      p10_bit_slice_6595 <= p10_data_enable ? p9_bit_slice_6595 : p10_bit_slice_6595;
      p10_bit_slice_6596 <= p10_data_enable ? p9_bit_slice_6596 : p10_bit_slice_6596;
      p10_bit_slice_6597 <= p10_data_enable ? p9_bit_slice_6597 : p10_bit_slice_6597;
      p10_bit_slice_6598 <= p10_data_enable ? p9_bit_slice_6598 : p10_bit_slice_6598;
      p10_bit_slice_6599 <= p10_data_enable ? p9_bit_slice_6599 : p10_bit_slice_6599;
      p10_bit_slice_6600 <= p10_data_enable ? p9_bit_slice_6600 : p10_bit_slice_6600;
      p10_bit_slice_6601 <= p10_data_enable ? p9_bit_slice_6601 : p10_bit_slice_6601;
      p10_bit_slice_6602 <= p10_data_enable ? p9_bit_slice_6602 : p10_bit_slice_6602;
      p10_bit_slice_6603 <= p10_data_enable ? p9_bit_slice_6603 : p10_bit_slice_6603;
      p10_bit_slice_6604 <= p10_data_enable ? p9_bit_slice_6604 : p10_bit_slice_6604;
      p10_bit_slice_6605 <= p10_data_enable ? p9_bit_slice_6605 : p10_bit_slice_6605;
      p10_bit_slice_6606 <= p10_data_enable ? p9_bit_slice_6606 : p10_bit_slice_6606;
      p10_bit_slice_6607 <= p10_data_enable ? p9_bit_slice_6607 : p10_bit_slice_6607;
      p10_negated <= p10_data_enable ? p9_negated : p10_negated;
      p11_b <= p11_data_enable ? p10_b : p11_b;
      p11_uge_6683 <= p11_data_enable ? p10_uge_6683 : p11_uge_6683;
      p11_bivisor__1 <= p11_data_enable ? p10_bivisor__1 : p11_bivisor__1;
      p11_uge_6691 <= p11_data_enable ? p10_uge_6691 : p11_uge_6691;
      p11_uge_6771 <= p11_data_enable ? p10_uge_6771 : p11_uge_6771;
      p11_uge_6851 <= p11_data_enable ? p10_uge_6851 : p11_uge_6851;
      p11_uge_6931 <= p11_data_enable ? p10_uge_6931 : p11_uge_6931;
      p11_uge_7011 <= p11_data_enable ? p10_uge_7011 : p11_uge_7011;
      p11_uge_7091 <= p11_data_enable ? p10_uge_7091 : p11_uge_7091;
      p11_uge_7171 <= p11_data_enable ? p10_uge_7171 : p11_uge_7171;
      p11_uge_7251 <= p11_data_enable ? p10_uge_7251 : p11_uge_7251;
      p11_uge_7331 <= p11_data_enable ? p10_uge_7331 : p11_uge_7331;
      p11_uge_7411 <= p11_data_enable ? p10_uge_7411 : p11_uge_7411;
      p11_concat_7490 <= p11_data_enable ? concat_7490 : p11_concat_7490;
      p11_uge_7491 <= p11_data_enable ? uge_7491 : p11_uge_7491;
      p11_bit_slice_6588 <= p11_data_enable ? p10_bit_slice_6588 : p11_bit_slice_6588;
      p11_bit_slice_6589 <= p11_data_enable ? p10_bit_slice_6589 : p11_bit_slice_6589;
      p11_bit_slice_6590 <= p11_data_enable ? p10_bit_slice_6590 : p11_bit_slice_6590;
      p11_bit_slice_6591 <= p11_data_enable ? p10_bit_slice_6591 : p11_bit_slice_6591;
      p11_bit_slice_6592 <= p11_data_enable ? p10_bit_slice_6592 : p11_bit_slice_6592;
      p11_bit_slice_6593 <= p11_data_enable ? p10_bit_slice_6593 : p11_bit_slice_6593;
      p11_bit_slice_6594 <= p11_data_enable ? p10_bit_slice_6594 : p11_bit_slice_6594;
      p11_bit_slice_6595 <= p11_data_enable ? p10_bit_slice_6595 : p11_bit_slice_6595;
      p11_bit_slice_6596 <= p11_data_enable ? p10_bit_slice_6596 : p11_bit_slice_6596;
      p11_bit_slice_6597 <= p11_data_enable ? p10_bit_slice_6597 : p11_bit_slice_6597;
      p11_bit_slice_6598 <= p11_data_enable ? p10_bit_slice_6598 : p11_bit_slice_6598;
      p11_bit_slice_6599 <= p11_data_enable ? p10_bit_slice_6599 : p11_bit_slice_6599;
      p11_bit_slice_6600 <= p11_data_enable ? p10_bit_slice_6600 : p11_bit_slice_6600;
      p11_bit_slice_6601 <= p11_data_enable ? p10_bit_slice_6601 : p11_bit_slice_6601;
      p11_bit_slice_6602 <= p11_data_enable ? p10_bit_slice_6602 : p11_bit_slice_6602;
      p11_bit_slice_6603 <= p11_data_enable ? p10_bit_slice_6603 : p11_bit_slice_6603;
      p11_bit_slice_6604 <= p11_data_enable ? p10_bit_slice_6604 : p11_bit_slice_6604;
      p11_bit_slice_6605 <= p11_data_enable ? p10_bit_slice_6605 : p11_bit_slice_6605;
      p11_bit_slice_6606 <= p11_data_enable ? p10_bit_slice_6606 : p11_bit_slice_6606;
      p11_bit_slice_6607 <= p11_data_enable ? p10_bit_slice_6607 : p11_bit_slice_6607;
      p11_negated <= p11_data_enable ? p10_negated : p11_negated;
      p12_b <= p12_data_enable ? p11_b : p12_b;
      p12_uge_6683 <= p12_data_enable ? p11_uge_6683 : p12_uge_6683;
      p12_bivisor__1 <= p12_data_enable ? p11_bivisor__1 : p12_bivisor__1;
      p12_uge_6691 <= p12_data_enable ? p11_uge_6691 : p12_uge_6691;
      p12_uge_6771 <= p12_data_enable ? p11_uge_6771 : p12_uge_6771;
      p12_uge_6851 <= p12_data_enable ? p11_uge_6851 : p12_uge_6851;
      p12_uge_6931 <= p12_data_enable ? p11_uge_6931 : p12_uge_6931;
      p12_uge_7011 <= p12_data_enable ? p11_uge_7011 : p12_uge_7011;
      p12_uge_7091 <= p12_data_enable ? p11_uge_7091 : p12_uge_7091;
      p12_uge_7171 <= p12_data_enable ? p11_uge_7171 : p12_uge_7171;
      p12_uge_7251 <= p12_data_enable ? p11_uge_7251 : p12_uge_7251;
      p12_uge_7331 <= p12_data_enable ? p11_uge_7331 : p12_uge_7331;
      p12_uge_7411 <= p12_data_enable ? p11_uge_7411 : p12_uge_7411;
      p12_uge_7491 <= p12_data_enable ? p11_uge_7491 : p12_uge_7491;
      p12_concat_7570 <= p12_data_enable ? concat_7570 : p12_concat_7570;
      p12_uge_7571 <= p12_data_enable ? uge_7571 : p12_uge_7571;
      p12_bit_slice_6589 <= p12_data_enable ? p11_bit_slice_6589 : p12_bit_slice_6589;
      p12_bit_slice_6590 <= p12_data_enable ? p11_bit_slice_6590 : p12_bit_slice_6590;
      p12_bit_slice_6591 <= p12_data_enable ? p11_bit_slice_6591 : p12_bit_slice_6591;
      p12_bit_slice_6592 <= p12_data_enable ? p11_bit_slice_6592 : p12_bit_slice_6592;
      p12_bit_slice_6593 <= p12_data_enable ? p11_bit_slice_6593 : p12_bit_slice_6593;
      p12_bit_slice_6594 <= p12_data_enable ? p11_bit_slice_6594 : p12_bit_slice_6594;
      p12_bit_slice_6595 <= p12_data_enable ? p11_bit_slice_6595 : p12_bit_slice_6595;
      p12_bit_slice_6596 <= p12_data_enable ? p11_bit_slice_6596 : p12_bit_slice_6596;
      p12_bit_slice_6597 <= p12_data_enable ? p11_bit_slice_6597 : p12_bit_slice_6597;
      p12_bit_slice_6598 <= p12_data_enable ? p11_bit_slice_6598 : p12_bit_slice_6598;
      p12_bit_slice_6599 <= p12_data_enable ? p11_bit_slice_6599 : p12_bit_slice_6599;
      p12_bit_slice_6600 <= p12_data_enable ? p11_bit_slice_6600 : p12_bit_slice_6600;
      p12_bit_slice_6601 <= p12_data_enable ? p11_bit_slice_6601 : p12_bit_slice_6601;
      p12_bit_slice_6602 <= p12_data_enable ? p11_bit_slice_6602 : p12_bit_slice_6602;
      p12_bit_slice_6603 <= p12_data_enable ? p11_bit_slice_6603 : p12_bit_slice_6603;
      p12_bit_slice_6604 <= p12_data_enable ? p11_bit_slice_6604 : p12_bit_slice_6604;
      p12_bit_slice_6605 <= p12_data_enable ? p11_bit_slice_6605 : p12_bit_slice_6605;
      p12_bit_slice_6606 <= p12_data_enable ? p11_bit_slice_6606 : p12_bit_slice_6606;
      p12_bit_slice_6607 <= p12_data_enable ? p11_bit_slice_6607 : p12_bit_slice_6607;
      p12_negated <= p12_data_enable ? p11_negated : p12_negated;
      p13_b <= p13_data_enable ? p12_b : p13_b;
      p13_uge_6683 <= p13_data_enable ? p12_uge_6683 : p13_uge_6683;
      p13_bivisor__1 <= p13_data_enable ? p12_bivisor__1 : p13_bivisor__1;
      p13_uge_6691 <= p13_data_enable ? p12_uge_6691 : p13_uge_6691;
      p13_uge_6771 <= p13_data_enable ? p12_uge_6771 : p13_uge_6771;
      p13_uge_6851 <= p13_data_enable ? p12_uge_6851 : p13_uge_6851;
      p13_uge_6931 <= p13_data_enable ? p12_uge_6931 : p13_uge_6931;
      p13_uge_7011 <= p13_data_enable ? p12_uge_7011 : p13_uge_7011;
      p13_uge_7091 <= p13_data_enable ? p12_uge_7091 : p13_uge_7091;
      p13_uge_7171 <= p13_data_enable ? p12_uge_7171 : p13_uge_7171;
      p13_uge_7251 <= p13_data_enable ? p12_uge_7251 : p13_uge_7251;
      p13_uge_7331 <= p13_data_enable ? p12_uge_7331 : p13_uge_7331;
      p13_uge_7411 <= p13_data_enable ? p12_uge_7411 : p13_uge_7411;
      p13_uge_7491 <= p13_data_enable ? p12_uge_7491 : p13_uge_7491;
      p13_uge_7571 <= p13_data_enable ? p12_uge_7571 : p13_uge_7571;
      p13_concat_7650 <= p13_data_enable ? concat_7650 : p13_concat_7650;
      p13_uge_7651 <= p13_data_enable ? uge_7651 : p13_uge_7651;
      p13_bit_slice_6590 <= p13_data_enable ? p12_bit_slice_6590 : p13_bit_slice_6590;
      p13_bit_slice_6591 <= p13_data_enable ? p12_bit_slice_6591 : p13_bit_slice_6591;
      p13_bit_slice_6592 <= p13_data_enable ? p12_bit_slice_6592 : p13_bit_slice_6592;
      p13_bit_slice_6593 <= p13_data_enable ? p12_bit_slice_6593 : p13_bit_slice_6593;
      p13_bit_slice_6594 <= p13_data_enable ? p12_bit_slice_6594 : p13_bit_slice_6594;
      p13_bit_slice_6595 <= p13_data_enable ? p12_bit_slice_6595 : p13_bit_slice_6595;
      p13_bit_slice_6596 <= p13_data_enable ? p12_bit_slice_6596 : p13_bit_slice_6596;
      p13_bit_slice_6597 <= p13_data_enable ? p12_bit_slice_6597 : p13_bit_slice_6597;
      p13_bit_slice_6598 <= p13_data_enable ? p12_bit_slice_6598 : p13_bit_slice_6598;
      p13_bit_slice_6599 <= p13_data_enable ? p12_bit_slice_6599 : p13_bit_slice_6599;
      p13_bit_slice_6600 <= p13_data_enable ? p12_bit_slice_6600 : p13_bit_slice_6600;
      p13_bit_slice_6601 <= p13_data_enable ? p12_bit_slice_6601 : p13_bit_slice_6601;
      p13_bit_slice_6602 <= p13_data_enable ? p12_bit_slice_6602 : p13_bit_slice_6602;
      p13_bit_slice_6603 <= p13_data_enable ? p12_bit_slice_6603 : p13_bit_slice_6603;
      p13_bit_slice_6604 <= p13_data_enable ? p12_bit_slice_6604 : p13_bit_slice_6604;
      p13_bit_slice_6605 <= p13_data_enable ? p12_bit_slice_6605 : p13_bit_slice_6605;
      p13_bit_slice_6606 <= p13_data_enable ? p12_bit_slice_6606 : p13_bit_slice_6606;
      p13_bit_slice_6607 <= p13_data_enable ? p12_bit_slice_6607 : p13_bit_slice_6607;
      p13_negated <= p13_data_enable ? p12_negated : p13_negated;
      p14_b <= p14_data_enable ? p13_b : p14_b;
      p14_uge_6683 <= p14_data_enable ? p13_uge_6683 : p14_uge_6683;
      p14_bivisor__1 <= p14_data_enable ? p13_bivisor__1 : p14_bivisor__1;
      p14_uge_6691 <= p14_data_enable ? p13_uge_6691 : p14_uge_6691;
      p14_uge_6771 <= p14_data_enable ? p13_uge_6771 : p14_uge_6771;
      p14_uge_6851 <= p14_data_enable ? p13_uge_6851 : p14_uge_6851;
      p14_uge_6931 <= p14_data_enable ? p13_uge_6931 : p14_uge_6931;
      p14_uge_7011 <= p14_data_enable ? p13_uge_7011 : p14_uge_7011;
      p14_uge_7091 <= p14_data_enable ? p13_uge_7091 : p14_uge_7091;
      p14_uge_7171 <= p14_data_enable ? p13_uge_7171 : p14_uge_7171;
      p14_uge_7251 <= p14_data_enable ? p13_uge_7251 : p14_uge_7251;
      p14_uge_7331 <= p14_data_enable ? p13_uge_7331 : p14_uge_7331;
      p14_uge_7411 <= p14_data_enable ? p13_uge_7411 : p14_uge_7411;
      p14_uge_7491 <= p14_data_enable ? p13_uge_7491 : p14_uge_7491;
      p14_uge_7571 <= p14_data_enable ? p13_uge_7571 : p14_uge_7571;
      p14_uge_7651 <= p14_data_enable ? p13_uge_7651 : p14_uge_7651;
      p14_concat_7730 <= p14_data_enable ? concat_7730 : p14_concat_7730;
      p14_uge_7731 <= p14_data_enable ? uge_7731 : p14_uge_7731;
      p14_bit_slice_6591 <= p14_data_enable ? p13_bit_slice_6591 : p14_bit_slice_6591;
      p14_bit_slice_6592 <= p14_data_enable ? p13_bit_slice_6592 : p14_bit_slice_6592;
      p14_bit_slice_6593 <= p14_data_enable ? p13_bit_slice_6593 : p14_bit_slice_6593;
      p14_bit_slice_6594 <= p14_data_enable ? p13_bit_slice_6594 : p14_bit_slice_6594;
      p14_bit_slice_6595 <= p14_data_enable ? p13_bit_slice_6595 : p14_bit_slice_6595;
      p14_bit_slice_6596 <= p14_data_enable ? p13_bit_slice_6596 : p14_bit_slice_6596;
      p14_bit_slice_6597 <= p14_data_enable ? p13_bit_slice_6597 : p14_bit_slice_6597;
      p14_bit_slice_6598 <= p14_data_enable ? p13_bit_slice_6598 : p14_bit_slice_6598;
      p14_bit_slice_6599 <= p14_data_enable ? p13_bit_slice_6599 : p14_bit_slice_6599;
      p14_bit_slice_6600 <= p14_data_enable ? p13_bit_slice_6600 : p14_bit_slice_6600;
      p14_bit_slice_6601 <= p14_data_enable ? p13_bit_slice_6601 : p14_bit_slice_6601;
      p14_bit_slice_6602 <= p14_data_enable ? p13_bit_slice_6602 : p14_bit_slice_6602;
      p14_bit_slice_6603 <= p14_data_enable ? p13_bit_slice_6603 : p14_bit_slice_6603;
      p14_bit_slice_6604 <= p14_data_enable ? p13_bit_slice_6604 : p14_bit_slice_6604;
      p14_bit_slice_6605 <= p14_data_enable ? p13_bit_slice_6605 : p14_bit_slice_6605;
      p14_bit_slice_6606 <= p14_data_enable ? p13_bit_slice_6606 : p14_bit_slice_6606;
      p14_bit_slice_6607 <= p14_data_enable ? p13_bit_slice_6607 : p14_bit_slice_6607;
      p14_negated <= p14_data_enable ? p13_negated : p14_negated;
      p15_b <= p15_data_enable ? p14_b : p15_b;
      p15_uge_6683 <= p15_data_enable ? p14_uge_6683 : p15_uge_6683;
      p15_bivisor__1 <= p15_data_enable ? p14_bivisor__1 : p15_bivisor__1;
      p15_uge_6691 <= p15_data_enable ? p14_uge_6691 : p15_uge_6691;
      p15_uge_6771 <= p15_data_enable ? p14_uge_6771 : p15_uge_6771;
      p15_uge_6851 <= p15_data_enable ? p14_uge_6851 : p15_uge_6851;
      p15_uge_6931 <= p15_data_enable ? p14_uge_6931 : p15_uge_6931;
      p15_uge_7011 <= p15_data_enable ? p14_uge_7011 : p15_uge_7011;
      p15_uge_7091 <= p15_data_enable ? p14_uge_7091 : p15_uge_7091;
      p15_uge_7171 <= p15_data_enable ? p14_uge_7171 : p15_uge_7171;
      p15_uge_7251 <= p15_data_enable ? p14_uge_7251 : p15_uge_7251;
      p15_uge_7331 <= p15_data_enable ? p14_uge_7331 : p15_uge_7331;
      p15_uge_7411 <= p15_data_enable ? p14_uge_7411 : p15_uge_7411;
      p15_uge_7491 <= p15_data_enable ? p14_uge_7491 : p15_uge_7491;
      p15_uge_7571 <= p15_data_enable ? p14_uge_7571 : p15_uge_7571;
      p15_uge_7651 <= p15_data_enable ? p14_uge_7651 : p15_uge_7651;
      p15_uge_7731 <= p15_data_enable ? p14_uge_7731 : p15_uge_7731;
      p15_concat_7810 <= p15_data_enable ? concat_7810 : p15_concat_7810;
      p15_uge_7811 <= p15_data_enable ? uge_7811 : p15_uge_7811;
      p15_bit_slice_6592 <= p15_data_enable ? p14_bit_slice_6592 : p15_bit_slice_6592;
      p15_bit_slice_6593 <= p15_data_enable ? p14_bit_slice_6593 : p15_bit_slice_6593;
      p15_bit_slice_6594 <= p15_data_enable ? p14_bit_slice_6594 : p15_bit_slice_6594;
      p15_bit_slice_6595 <= p15_data_enable ? p14_bit_slice_6595 : p15_bit_slice_6595;
      p15_bit_slice_6596 <= p15_data_enable ? p14_bit_slice_6596 : p15_bit_slice_6596;
      p15_bit_slice_6597 <= p15_data_enable ? p14_bit_slice_6597 : p15_bit_slice_6597;
      p15_bit_slice_6598 <= p15_data_enable ? p14_bit_slice_6598 : p15_bit_slice_6598;
      p15_bit_slice_6599 <= p15_data_enable ? p14_bit_slice_6599 : p15_bit_slice_6599;
      p15_bit_slice_6600 <= p15_data_enable ? p14_bit_slice_6600 : p15_bit_slice_6600;
      p15_bit_slice_6601 <= p15_data_enable ? p14_bit_slice_6601 : p15_bit_slice_6601;
      p15_bit_slice_6602 <= p15_data_enable ? p14_bit_slice_6602 : p15_bit_slice_6602;
      p15_bit_slice_6603 <= p15_data_enable ? p14_bit_slice_6603 : p15_bit_slice_6603;
      p15_bit_slice_6604 <= p15_data_enable ? p14_bit_slice_6604 : p15_bit_slice_6604;
      p15_bit_slice_6605 <= p15_data_enable ? p14_bit_slice_6605 : p15_bit_slice_6605;
      p15_bit_slice_6606 <= p15_data_enable ? p14_bit_slice_6606 : p15_bit_slice_6606;
      p15_bit_slice_6607 <= p15_data_enable ? p14_bit_slice_6607 : p15_bit_slice_6607;
      p15_negated <= p15_data_enable ? p14_negated : p15_negated;
      p16_b <= p16_data_enable ? p15_b : p16_b;
      p16_uge_6683 <= p16_data_enable ? p15_uge_6683 : p16_uge_6683;
      p16_bivisor__1 <= p16_data_enable ? p15_bivisor__1 : p16_bivisor__1;
      p16_uge_6691 <= p16_data_enable ? p15_uge_6691 : p16_uge_6691;
      p16_uge_6771 <= p16_data_enable ? p15_uge_6771 : p16_uge_6771;
      p16_uge_6851 <= p16_data_enable ? p15_uge_6851 : p16_uge_6851;
      p16_uge_6931 <= p16_data_enable ? p15_uge_6931 : p16_uge_6931;
      p16_uge_7011 <= p16_data_enable ? p15_uge_7011 : p16_uge_7011;
      p16_uge_7091 <= p16_data_enable ? p15_uge_7091 : p16_uge_7091;
      p16_uge_7171 <= p16_data_enable ? p15_uge_7171 : p16_uge_7171;
      p16_uge_7251 <= p16_data_enable ? p15_uge_7251 : p16_uge_7251;
      p16_uge_7331 <= p16_data_enable ? p15_uge_7331 : p16_uge_7331;
      p16_uge_7411 <= p16_data_enable ? p15_uge_7411 : p16_uge_7411;
      p16_uge_7491 <= p16_data_enable ? p15_uge_7491 : p16_uge_7491;
      p16_uge_7571 <= p16_data_enable ? p15_uge_7571 : p16_uge_7571;
      p16_uge_7651 <= p16_data_enable ? p15_uge_7651 : p16_uge_7651;
      p16_uge_7731 <= p16_data_enable ? p15_uge_7731 : p16_uge_7731;
      p16_uge_7811 <= p16_data_enable ? p15_uge_7811 : p16_uge_7811;
      p16_concat_7890 <= p16_data_enable ? concat_7890 : p16_concat_7890;
      p16_uge_7891 <= p16_data_enable ? uge_7891 : p16_uge_7891;
      p16_bit_slice_6593 <= p16_data_enable ? p15_bit_slice_6593 : p16_bit_slice_6593;
      p16_bit_slice_6594 <= p16_data_enable ? p15_bit_slice_6594 : p16_bit_slice_6594;
      p16_bit_slice_6595 <= p16_data_enable ? p15_bit_slice_6595 : p16_bit_slice_6595;
      p16_bit_slice_6596 <= p16_data_enable ? p15_bit_slice_6596 : p16_bit_slice_6596;
      p16_bit_slice_6597 <= p16_data_enable ? p15_bit_slice_6597 : p16_bit_slice_6597;
      p16_bit_slice_6598 <= p16_data_enable ? p15_bit_slice_6598 : p16_bit_slice_6598;
      p16_bit_slice_6599 <= p16_data_enable ? p15_bit_slice_6599 : p16_bit_slice_6599;
      p16_bit_slice_6600 <= p16_data_enable ? p15_bit_slice_6600 : p16_bit_slice_6600;
      p16_bit_slice_6601 <= p16_data_enable ? p15_bit_slice_6601 : p16_bit_slice_6601;
      p16_bit_slice_6602 <= p16_data_enable ? p15_bit_slice_6602 : p16_bit_slice_6602;
      p16_bit_slice_6603 <= p16_data_enable ? p15_bit_slice_6603 : p16_bit_slice_6603;
      p16_bit_slice_6604 <= p16_data_enable ? p15_bit_slice_6604 : p16_bit_slice_6604;
      p16_bit_slice_6605 <= p16_data_enable ? p15_bit_slice_6605 : p16_bit_slice_6605;
      p16_bit_slice_6606 <= p16_data_enable ? p15_bit_slice_6606 : p16_bit_slice_6606;
      p16_bit_slice_6607 <= p16_data_enable ? p15_bit_slice_6607 : p16_bit_slice_6607;
      p16_negated <= p16_data_enable ? p15_negated : p16_negated;
      p17_b <= p17_data_enable ? p16_b : p17_b;
      p17_uge_6683 <= p17_data_enable ? p16_uge_6683 : p17_uge_6683;
      p17_bivisor__1 <= p17_data_enable ? p16_bivisor__1 : p17_bivisor__1;
      p17_uge_6691 <= p17_data_enable ? p16_uge_6691 : p17_uge_6691;
      p17_uge_6771 <= p17_data_enable ? p16_uge_6771 : p17_uge_6771;
      p17_uge_6851 <= p17_data_enable ? p16_uge_6851 : p17_uge_6851;
      p17_uge_6931 <= p17_data_enable ? p16_uge_6931 : p17_uge_6931;
      p17_uge_7011 <= p17_data_enable ? p16_uge_7011 : p17_uge_7011;
      p17_uge_7091 <= p17_data_enable ? p16_uge_7091 : p17_uge_7091;
      p17_uge_7171 <= p17_data_enable ? p16_uge_7171 : p17_uge_7171;
      p17_uge_7251 <= p17_data_enable ? p16_uge_7251 : p17_uge_7251;
      p17_uge_7331 <= p17_data_enable ? p16_uge_7331 : p17_uge_7331;
      p17_uge_7411 <= p17_data_enable ? p16_uge_7411 : p17_uge_7411;
      p17_uge_7491 <= p17_data_enable ? p16_uge_7491 : p17_uge_7491;
      p17_uge_7571 <= p17_data_enable ? p16_uge_7571 : p17_uge_7571;
      p17_uge_7651 <= p17_data_enable ? p16_uge_7651 : p17_uge_7651;
      p17_uge_7731 <= p17_data_enable ? p16_uge_7731 : p17_uge_7731;
      p17_uge_7811 <= p17_data_enable ? p16_uge_7811 : p17_uge_7811;
      p17_uge_7891 <= p17_data_enable ? p16_uge_7891 : p17_uge_7891;
      p17_concat_7970 <= p17_data_enable ? concat_7970 : p17_concat_7970;
      p17_uge_7971 <= p17_data_enable ? uge_7971 : p17_uge_7971;
      p17_bit_slice_6594 <= p17_data_enable ? p16_bit_slice_6594 : p17_bit_slice_6594;
      p17_bit_slice_6595 <= p17_data_enable ? p16_bit_slice_6595 : p17_bit_slice_6595;
      p17_bit_slice_6596 <= p17_data_enable ? p16_bit_slice_6596 : p17_bit_slice_6596;
      p17_bit_slice_6597 <= p17_data_enable ? p16_bit_slice_6597 : p17_bit_slice_6597;
      p17_bit_slice_6598 <= p17_data_enable ? p16_bit_slice_6598 : p17_bit_slice_6598;
      p17_bit_slice_6599 <= p17_data_enable ? p16_bit_slice_6599 : p17_bit_slice_6599;
      p17_bit_slice_6600 <= p17_data_enable ? p16_bit_slice_6600 : p17_bit_slice_6600;
      p17_bit_slice_6601 <= p17_data_enable ? p16_bit_slice_6601 : p17_bit_slice_6601;
      p17_bit_slice_6602 <= p17_data_enable ? p16_bit_slice_6602 : p17_bit_slice_6602;
      p17_bit_slice_6603 <= p17_data_enable ? p16_bit_slice_6603 : p17_bit_slice_6603;
      p17_bit_slice_6604 <= p17_data_enable ? p16_bit_slice_6604 : p17_bit_slice_6604;
      p17_bit_slice_6605 <= p17_data_enable ? p16_bit_slice_6605 : p17_bit_slice_6605;
      p17_bit_slice_6606 <= p17_data_enable ? p16_bit_slice_6606 : p17_bit_slice_6606;
      p17_bit_slice_6607 <= p17_data_enable ? p16_bit_slice_6607 : p17_bit_slice_6607;
      p17_negated <= p17_data_enable ? p16_negated : p17_negated;
      p18_b <= p18_data_enable ? p17_b : p18_b;
      p18_uge_6683 <= p18_data_enable ? p17_uge_6683 : p18_uge_6683;
      p18_bivisor__1 <= p18_data_enable ? p17_bivisor__1 : p18_bivisor__1;
      p18_uge_6691 <= p18_data_enable ? p17_uge_6691 : p18_uge_6691;
      p18_uge_6771 <= p18_data_enable ? p17_uge_6771 : p18_uge_6771;
      p18_uge_6851 <= p18_data_enable ? p17_uge_6851 : p18_uge_6851;
      p18_uge_6931 <= p18_data_enable ? p17_uge_6931 : p18_uge_6931;
      p18_uge_7011 <= p18_data_enable ? p17_uge_7011 : p18_uge_7011;
      p18_uge_7091 <= p18_data_enable ? p17_uge_7091 : p18_uge_7091;
      p18_uge_7171 <= p18_data_enable ? p17_uge_7171 : p18_uge_7171;
      p18_uge_7251 <= p18_data_enable ? p17_uge_7251 : p18_uge_7251;
      p18_uge_7331 <= p18_data_enable ? p17_uge_7331 : p18_uge_7331;
      p18_uge_7411 <= p18_data_enable ? p17_uge_7411 : p18_uge_7411;
      p18_uge_7491 <= p18_data_enable ? p17_uge_7491 : p18_uge_7491;
      p18_uge_7571 <= p18_data_enable ? p17_uge_7571 : p18_uge_7571;
      p18_uge_7651 <= p18_data_enable ? p17_uge_7651 : p18_uge_7651;
      p18_uge_7731 <= p18_data_enable ? p17_uge_7731 : p18_uge_7731;
      p18_uge_7811 <= p18_data_enable ? p17_uge_7811 : p18_uge_7811;
      p18_uge_7891 <= p18_data_enable ? p17_uge_7891 : p18_uge_7891;
      p18_uge_7971 <= p18_data_enable ? p17_uge_7971 : p18_uge_7971;
      p18_concat_8050 <= p18_data_enable ? concat_8050 : p18_concat_8050;
      p18_uge_8051 <= p18_data_enable ? uge_8051 : p18_uge_8051;
      p18_bit_slice_6595 <= p18_data_enable ? p17_bit_slice_6595 : p18_bit_slice_6595;
      p18_bit_slice_6596 <= p18_data_enable ? p17_bit_slice_6596 : p18_bit_slice_6596;
      p18_bit_slice_6597 <= p18_data_enable ? p17_bit_slice_6597 : p18_bit_slice_6597;
      p18_bit_slice_6598 <= p18_data_enable ? p17_bit_slice_6598 : p18_bit_slice_6598;
      p18_bit_slice_6599 <= p18_data_enable ? p17_bit_slice_6599 : p18_bit_slice_6599;
      p18_bit_slice_6600 <= p18_data_enable ? p17_bit_slice_6600 : p18_bit_slice_6600;
      p18_bit_slice_6601 <= p18_data_enable ? p17_bit_slice_6601 : p18_bit_slice_6601;
      p18_bit_slice_6602 <= p18_data_enable ? p17_bit_slice_6602 : p18_bit_slice_6602;
      p18_bit_slice_6603 <= p18_data_enable ? p17_bit_slice_6603 : p18_bit_slice_6603;
      p18_bit_slice_6604 <= p18_data_enable ? p17_bit_slice_6604 : p18_bit_slice_6604;
      p18_bit_slice_6605 <= p18_data_enable ? p17_bit_slice_6605 : p18_bit_slice_6605;
      p18_bit_slice_6606 <= p18_data_enable ? p17_bit_slice_6606 : p18_bit_slice_6606;
      p18_bit_slice_6607 <= p18_data_enable ? p17_bit_slice_6607 : p18_bit_slice_6607;
      p18_negated <= p18_data_enable ? p17_negated : p18_negated;
      p19_b <= p19_data_enable ? p18_b : p19_b;
      p19_uge_6683 <= p19_data_enable ? p18_uge_6683 : p19_uge_6683;
      p19_bivisor__1 <= p19_data_enable ? p18_bivisor__1 : p19_bivisor__1;
      p19_uge_6691 <= p19_data_enable ? p18_uge_6691 : p19_uge_6691;
      p19_uge_6771 <= p19_data_enable ? p18_uge_6771 : p19_uge_6771;
      p19_uge_6851 <= p19_data_enable ? p18_uge_6851 : p19_uge_6851;
      p19_uge_6931 <= p19_data_enable ? p18_uge_6931 : p19_uge_6931;
      p19_uge_7011 <= p19_data_enable ? p18_uge_7011 : p19_uge_7011;
      p19_uge_7091 <= p19_data_enable ? p18_uge_7091 : p19_uge_7091;
      p19_uge_7171 <= p19_data_enable ? p18_uge_7171 : p19_uge_7171;
      p19_uge_7251 <= p19_data_enable ? p18_uge_7251 : p19_uge_7251;
      p19_uge_7331 <= p19_data_enable ? p18_uge_7331 : p19_uge_7331;
      p19_uge_7411 <= p19_data_enable ? p18_uge_7411 : p19_uge_7411;
      p19_uge_7491 <= p19_data_enable ? p18_uge_7491 : p19_uge_7491;
      p19_uge_7571 <= p19_data_enable ? p18_uge_7571 : p19_uge_7571;
      p19_uge_7651 <= p19_data_enable ? p18_uge_7651 : p19_uge_7651;
      p19_uge_7731 <= p19_data_enable ? p18_uge_7731 : p19_uge_7731;
      p19_uge_7811 <= p19_data_enable ? p18_uge_7811 : p19_uge_7811;
      p19_uge_7891 <= p19_data_enable ? p18_uge_7891 : p19_uge_7891;
      p19_uge_7971 <= p19_data_enable ? p18_uge_7971 : p19_uge_7971;
      p19_uge_8051 <= p19_data_enable ? p18_uge_8051 : p19_uge_8051;
      p19_concat_8130 <= p19_data_enable ? concat_8130 : p19_concat_8130;
      p19_uge_8131 <= p19_data_enable ? uge_8131 : p19_uge_8131;
      p19_bit_slice_6596 <= p19_data_enable ? p18_bit_slice_6596 : p19_bit_slice_6596;
      p19_bit_slice_6597 <= p19_data_enable ? p18_bit_slice_6597 : p19_bit_slice_6597;
      p19_bit_slice_6598 <= p19_data_enable ? p18_bit_slice_6598 : p19_bit_slice_6598;
      p19_bit_slice_6599 <= p19_data_enable ? p18_bit_slice_6599 : p19_bit_slice_6599;
      p19_bit_slice_6600 <= p19_data_enable ? p18_bit_slice_6600 : p19_bit_slice_6600;
      p19_bit_slice_6601 <= p19_data_enable ? p18_bit_slice_6601 : p19_bit_slice_6601;
      p19_bit_slice_6602 <= p19_data_enable ? p18_bit_slice_6602 : p19_bit_slice_6602;
      p19_bit_slice_6603 <= p19_data_enable ? p18_bit_slice_6603 : p19_bit_slice_6603;
      p19_bit_slice_6604 <= p19_data_enable ? p18_bit_slice_6604 : p19_bit_slice_6604;
      p19_bit_slice_6605 <= p19_data_enable ? p18_bit_slice_6605 : p19_bit_slice_6605;
      p19_bit_slice_6606 <= p19_data_enable ? p18_bit_slice_6606 : p19_bit_slice_6606;
      p19_bit_slice_6607 <= p19_data_enable ? p18_bit_slice_6607 : p19_bit_slice_6607;
      p19_negated <= p19_data_enable ? p18_negated : p19_negated;
      p20_b <= p20_data_enable ? p19_b : p20_b;
      p20_uge_6683 <= p20_data_enable ? p19_uge_6683 : p20_uge_6683;
      p20_bivisor__1 <= p20_data_enable ? p19_bivisor__1 : p20_bivisor__1;
      p20_uge_6691 <= p20_data_enable ? p19_uge_6691 : p20_uge_6691;
      p20_uge_6771 <= p20_data_enable ? p19_uge_6771 : p20_uge_6771;
      p20_uge_6851 <= p20_data_enable ? p19_uge_6851 : p20_uge_6851;
      p20_uge_6931 <= p20_data_enable ? p19_uge_6931 : p20_uge_6931;
      p20_uge_7011 <= p20_data_enable ? p19_uge_7011 : p20_uge_7011;
      p20_uge_7091 <= p20_data_enable ? p19_uge_7091 : p20_uge_7091;
      p20_uge_7171 <= p20_data_enable ? p19_uge_7171 : p20_uge_7171;
      p20_uge_7251 <= p20_data_enable ? p19_uge_7251 : p20_uge_7251;
      p20_uge_7331 <= p20_data_enable ? p19_uge_7331 : p20_uge_7331;
      p20_uge_7411 <= p20_data_enable ? p19_uge_7411 : p20_uge_7411;
      p20_uge_7491 <= p20_data_enable ? p19_uge_7491 : p20_uge_7491;
      p20_uge_7571 <= p20_data_enable ? p19_uge_7571 : p20_uge_7571;
      p20_uge_7651 <= p20_data_enable ? p19_uge_7651 : p20_uge_7651;
      p20_uge_7731 <= p20_data_enable ? p19_uge_7731 : p20_uge_7731;
      p20_uge_7811 <= p20_data_enable ? p19_uge_7811 : p20_uge_7811;
      p20_uge_7891 <= p20_data_enable ? p19_uge_7891 : p20_uge_7891;
      p20_uge_7971 <= p20_data_enable ? p19_uge_7971 : p20_uge_7971;
      p20_uge_8051 <= p20_data_enable ? p19_uge_8051 : p20_uge_8051;
      p20_uge_8131 <= p20_data_enable ? p19_uge_8131 : p20_uge_8131;
      p20_concat_8210 <= p20_data_enable ? concat_8210 : p20_concat_8210;
      p20_uge_8211 <= p20_data_enable ? uge_8211 : p20_uge_8211;
      p20_bit_slice_6597 <= p20_data_enable ? p19_bit_slice_6597 : p20_bit_slice_6597;
      p20_bit_slice_6598 <= p20_data_enable ? p19_bit_slice_6598 : p20_bit_slice_6598;
      p20_bit_slice_6599 <= p20_data_enable ? p19_bit_slice_6599 : p20_bit_slice_6599;
      p20_bit_slice_6600 <= p20_data_enable ? p19_bit_slice_6600 : p20_bit_slice_6600;
      p20_bit_slice_6601 <= p20_data_enable ? p19_bit_slice_6601 : p20_bit_slice_6601;
      p20_bit_slice_6602 <= p20_data_enable ? p19_bit_slice_6602 : p20_bit_slice_6602;
      p20_bit_slice_6603 <= p20_data_enable ? p19_bit_slice_6603 : p20_bit_slice_6603;
      p20_bit_slice_6604 <= p20_data_enable ? p19_bit_slice_6604 : p20_bit_slice_6604;
      p20_bit_slice_6605 <= p20_data_enable ? p19_bit_slice_6605 : p20_bit_slice_6605;
      p20_bit_slice_6606 <= p20_data_enable ? p19_bit_slice_6606 : p20_bit_slice_6606;
      p20_bit_slice_6607 <= p20_data_enable ? p19_bit_slice_6607 : p20_bit_slice_6607;
      p20_negated <= p20_data_enable ? p19_negated : p20_negated;
      p21_b <= p21_data_enable ? p20_b : p21_b;
      p21_uge_6683 <= p21_data_enable ? p20_uge_6683 : p21_uge_6683;
      p21_bivisor__1 <= p21_data_enable ? p20_bivisor__1 : p21_bivisor__1;
      p21_uge_6691 <= p21_data_enable ? p20_uge_6691 : p21_uge_6691;
      p21_uge_6771 <= p21_data_enable ? p20_uge_6771 : p21_uge_6771;
      p21_uge_6851 <= p21_data_enable ? p20_uge_6851 : p21_uge_6851;
      p21_uge_6931 <= p21_data_enable ? p20_uge_6931 : p21_uge_6931;
      p21_uge_7011 <= p21_data_enable ? p20_uge_7011 : p21_uge_7011;
      p21_uge_7091 <= p21_data_enable ? p20_uge_7091 : p21_uge_7091;
      p21_uge_7171 <= p21_data_enable ? p20_uge_7171 : p21_uge_7171;
      p21_uge_7251 <= p21_data_enable ? p20_uge_7251 : p21_uge_7251;
      p21_uge_7331 <= p21_data_enable ? p20_uge_7331 : p21_uge_7331;
      p21_uge_7411 <= p21_data_enable ? p20_uge_7411 : p21_uge_7411;
      p21_uge_7491 <= p21_data_enable ? p20_uge_7491 : p21_uge_7491;
      p21_uge_7571 <= p21_data_enable ? p20_uge_7571 : p21_uge_7571;
      p21_uge_7651 <= p21_data_enable ? p20_uge_7651 : p21_uge_7651;
      p21_uge_7731 <= p21_data_enable ? p20_uge_7731 : p21_uge_7731;
      p21_uge_7811 <= p21_data_enable ? p20_uge_7811 : p21_uge_7811;
      p21_uge_7891 <= p21_data_enable ? p20_uge_7891 : p21_uge_7891;
      p21_uge_7971 <= p21_data_enable ? p20_uge_7971 : p21_uge_7971;
      p21_uge_8051 <= p21_data_enable ? p20_uge_8051 : p21_uge_8051;
      p21_uge_8131 <= p21_data_enable ? p20_uge_8131 : p21_uge_8131;
      p21_uge_8211 <= p21_data_enable ? p20_uge_8211 : p21_uge_8211;
      p21_concat_8290 <= p21_data_enable ? concat_8290 : p21_concat_8290;
      p21_uge_8291 <= p21_data_enable ? uge_8291 : p21_uge_8291;
      p21_bit_slice_6598 <= p21_data_enable ? p20_bit_slice_6598 : p21_bit_slice_6598;
      p21_bit_slice_6599 <= p21_data_enable ? p20_bit_slice_6599 : p21_bit_slice_6599;
      p21_bit_slice_6600 <= p21_data_enable ? p20_bit_slice_6600 : p21_bit_slice_6600;
      p21_bit_slice_6601 <= p21_data_enable ? p20_bit_slice_6601 : p21_bit_slice_6601;
      p21_bit_slice_6602 <= p21_data_enable ? p20_bit_slice_6602 : p21_bit_slice_6602;
      p21_bit_slice_6603 <= p21_data_enable ? p20_bit_slice_6603 : p21_bit_slice_6603;
      p21_bit_slice_6604 <= p21_data_enable ? p20_bit_slice_6604 : p21_bit_slice_6604;
      p21_bit_slice_6605 <= p21_data_enable ? p20_bit_slice_6605 : p21_bit_slice_6605;
      p21_bit_slice_6606 <= p21_data_enable ? p20_bit_slice_6606 : p21_bit_slice_6606;
      p21_bit_slice_6607 <= p21_data_enable ? p20_bit_slice_6607 : p21_bit_slice_6607;
      p21_negated <= p21_data_enable ? p20_negated : p21_negated;
      p22_b <= p22_data_enable ? p21_b : p22_b;
      p22_uge_6683 <= p22_data_enable ? p21_uge_6683 : p22_uge_6683;
      p22_bivisor__1 <= p22_data_enable ? p21_bivisor__1 : p22_bivisor__1;
      p22_uge_6691 <= p22_data_enable ? p21_uge_6691 : p22_uge_6691;
      p22_uge_6771 <= p22_data_enable ? p21_uge_6771 : p22_uge_6771;
      p22_uge_6851 <= p22_data_enable ? p21_uge_6851 : p22_uge_6851;
      p22_uge_6931 <= p22_data_enable ? p21_uge_6931 : p22_uge_6931;
      p22_uge_7011 <= p22_data_enable ? p21_uge_7011 : p22_uge_7011;
      p22_uge_7091 <= p22_data_enable ? p21_uge_7091 : p22_uge_7091;
      p22_uge_7171 <= p22_data_enable ? p21_uge_7171 : p22_uge_7171;
      p22_uge_7251 <= p22_data_enable ? p21_uge_7251 : p22_uge_7251;
      p22_uge_7331 <= p22_data_enable ? p21_uge_7331 : p22_uge_7331;
      p22_uge_7411 <= p22_data_enable ? p21_uge_7411 : p22_uge_7411;
      p22_uge_7491 <= p22_data_enable ? p21_uge_7491 : p22_uge_7491;
      p22_uge_7571 <= p22_data_enable ? p21_uge_7571 : p22_uge_7571;
      p22_uge_7651 <= p22_data_enable ? p21_uge_7651 : p22_uge_7651;
      p22_uge_7731 <= p22_data_enable ? p21_uge_7731 : p22_uge_7731;
      p22_uge_7811 <= p22_data_enable ? p21_uge_7811 : p22_uge_7811;
      p22_uge_7891 <= p22_data_enable ? p21_uge_7891 : p22_uge_7891;
      p22_uge_7971 <= p22_data_enable ? p21_uge_7971 : p22_uge_7971;
      p22_uge_8051 <= p22_data_enable ? p21_uge_8051 : p22_uge_8051;
      p22_uge_8131 <= p22_data_enable ? p21_uge_8131 : p22_uge_8131;
      p22_uge_8211 <= p22_data_enable ? p21_uge_8211 : p22_uge_8211;
      p22_uge_8291 <= p22_data_enable ? p21_uge_8291 : p22_uge_8291;
      p22_concat_8370 <= p22_data_enable ? concat_8370 : p22_concat_8370;
      p22_uge_8371 <= p22_data_enable ? uge_8371 : p22_uge_8371;
      p22_bit_slice_6599 <= p22_data_enable ? p21_bit_slice_6599 : p22_bit_slice_6599;
      p22_bit_slice_6600 <= p22_data_enable ? p21_bit_slice_6600 : p22_bit_slice_6600;
      p22_bit_slice_6601 <= p22_data_enable ? p21_bit_slice_6601 : p22_bit_slice_6601;
      p22_bit_slice_6602 <= p22_data_enable ? p21_bit_slice_6602 : p22_bit_slice_6602;
      p22_bit_slice_6603 <= p22_data_enable ? p21_bit_slice_6603 : p22_bit_slice_6603;
      p22_bit_slice_6604 <= p22_data_enable ? p21_bit_slice_6604 : p22_bit_slice_6604;
      p22_bit_slice_6605 <= p22_data_enable ? p21_bit_slice_6605 : p22_bit_slice_6605;
      p22_bit_slice_6606 <= p22_data_enable ? p21_bit_slice_6606 : p22_bit_slice_6606;
      p22_bit_slice_6607 <= p22_data_enable ? p21_bit_slice_6607 : p22_bit_slice_6607;
      p22_negated <= p22_data_enable ? p21_negated : p22_negated;
      p23_b <= p23_data_enable ? p22_b : p23_b;
      p23_uge_6683 <= p23_data_enable ? p22_uge_6683 : p23_uge_6683;
      p23_bivisor__1 <= p23_data_enable ? p22_bivisor__1 : p23_bivisor__1;
      p23_uge_6691 <= p23_data_enable ? p22_uge_6691 : p23_uge_6691;
      p23_uge_6771 <= p23_data_enable ? p22_uge_6771 : p23_uge_6771;
      p23_uge_6851 <= p23_data_enable ? p22_uge_6851 : p23_uge_6851;
      p23_uge_6931 <= p23_data_enable ? p22_uge_6931 : p23_uge_6931;
      p23_uge_7011 <= p23_data_enable ? p22_uge_7011 : p23_uge_7011;
      p23_uge_7091 <= p23_data_enable ? p22_uge_7091 : p23_uge_7091;
      p23_uge_7171 <= p23_data_enable ? p22_uge_7171 : p23_uge_7171;
      p23_uge_7251 <= p23_data_enable ? p22_uge_7251 : p23_uge_7251;
      p23_uge_7331 <= p23_data_enable ? p22_uge_7331 : p23_uge_7331;
      p23_uge_7411 <= p23_data_enable ? p22_uge_7411 : p23_uge_7411;
      p23_uge_7491 <= p23_data_enable ? p22_uge_7491 : p23_uge_7491;
      p23_uge_7571 <= p23_data_enable ? p22_uge_7571 : p23_uge_7571;
      p23_uge_7651 <= p23_data_enable ? p22_uge_7651 : p23_uge_7651;
      p23_uge_7731 <= p23_data_enable ? p22_uge_7731 : p23_uge_7731;
      p23_uge_7811 <= p23_data_enable ? p22_uge_7811 : p23_uge_7811;
      p23_uge_7891 <= p23_data_enable ? p22_uge_7891 : p23_uge_7891;
      p23_uge_7971 <= p23_data_enable ? p22_uge_7971 : p23_uge_7971;
      p23_uge_8051 <= p23_data_enable ? p22_uge_8051 : p23_uge_8051;
      p23_uge_8131 <= p23_data_enable ? p22_uge_8131 : p23_uge_8131;
      p23_uge_8211 <= p23_data_enable ? p22_uge_8211 : p23_uge_8211;
      p23_uge_8291 <= p23_data_enable ? p22_uge_8291 : p23_uge_8291;
      p23_uge_8371 <= p23_data_enable ? p22_uge_8371 : p23_uge_8371;
      p23_concat_8450 <= p23_data_enable ? concat_8450 : p23_concat_8450;
      p23_uge_8451 <= p23_data_enable ? uge_8451 : p23_uge_8451;
      p23_bit_slice_6600 <= p23_data_enable ? p22_bit_slice_6600 : p23_bit_slice_6600;
      p23_bit_slice_6601 <= p23_data_enable ? p22_bit_slice_6601 : p23_bit_slice_6601;
      p23_bit_slice_6602 <= p23_data_enable ? p22_bit_slice_6602 : p23_bit_slice_6602;
      p23_bit_slice_6603 <= p23_data_enable ? p22_bit_slice_6603 : p23_bit_slice_6603;
      p23_bit_slice_6604 <= p23_data_enable ? p22_bit_slice_6604 : p23_bit_slice_6604;
      p23_bit_slice_6605 <= p23_data_enable ? p22_bit_slice_6605 : p23_bit_slice_6605;
      p23_bit_slice_6606 <= p23_data_enable ? p22_bit_slice_6606 : p23_bit_slice_6606;
      p23_bit_slice_6607 <= p23_data_enable ? p22_bit_slice_6607 : p23_bit_slice_6607;
      p23_negated <= p23_data_enable ? p22_negated : p23_negated;
      p24_b <= p24_data_enable ? p23_b : p24_b;
      p24_uge_6683 <= p24_data_enable ? p23_uge_6683 : p24_uge_6683;
      p24_bivisor__1 <= p24_data_enable ? p23_bivisor__1 : p24_bivisor__1;
      p24_uge_6691 <= p24_data_enable ? p23_uge_6691 : p24_uge_6691;
      p24_uge_6771 <= p24_data_enable ? p23_uge_6771 : p24_uge_6771;
      p24_uge_6851 <= p24_data_enable ? p23_uge_6851 : p24_uge_6851;
      p24_uge_6931 <= p24_data_enable ? p23_uge_6931 : p24_uge_6931;
      p24_uge_7011 <= p24_data_enable ? p23_uge_7011 : p24_uge_7011;
      p24_uge_7091 <= p24_data_enable ? p23_uge_7091 : p24_uge_7091;
      p24_uge_7171 <= p24_data_enable ? p23_uge_7171 : p24_uge_7171;
      p24_uge_7251 <= p24_data_enable ? p23_uge_7251 : p24_uge_7251;
      p24_uge_7331 <= p24_data_enable ? p23_uge_7331 : p24_uge_7331;
      p24_uge_7411 <= p24_data_enable ? p23_uge_7411 : p24_uge_7411;
      p24_uge_7491 <= p24_data_enable ? p23_uge_7491 : p24_uge_7491;
      p24_uge_7571 <= p24_data_enable ? p23_uge_7571 : p24_uge_7571;
      p24_uge_7651 <= p24_data_enable ? p23_uge_7651 : p24_uge_7651;
      p24_uge_7731 <= p24_data_enable ? p23_uge_7731 : p24_uge_7731;
      p24_uge_7811 <= p24_data_enable ? p23_uge_7811 : p24_uge_7811;
      p24_uge_7891 <= p24_data_enable ? p23_uge_7891 : p24_uge_7891;
      p24_uge_7971 <= p24_data_enable ? p23_uge_7971 : p24_uge_7971;
      p24_uge_8051 <= p24_data_enable ? p23_uge_8051 : p24_uge_8051;
      p24_uge_8131 <= p24_data_enable ? p23_uge_8131 : p24_uge_8131;
      p24_uge_8211 <= p24_data_enable ? p23_uge_8211 : p24_uge_8211;
      p24_uge_8291 <= p24_data_enable ? p23_uge_8291 : p24_uge_8291;
      p24_uge_8371 <= p24_data_enable ? p23_uge_8371 : p24_uge_8371;
      p24_uge_8451 <= p24_data_enable ? p23_uge_8451 : p24_uge_8451;
      p24_concat_8530 <= p24_data_enable ? concat_8530 : p24_concat_8530;
      p24_uge_8531 <= p24_data_enable ? uge_8531 : p24_uge_8531;
      p24_bit_slice_6601 <= p24_data_enable ? p23_bit_slice_6601 : p24_bit_slice_6601;
      p24_bit_slice_6602 <= p24_data_enable ? p23_bit_slice_6602 : p24_bit_slice_6602;
      p24_bit_slice_6603 <= p24_data_enable ? p23_bit_slice_6603 : p24_bit_slice_6603;
      p24_bit_slice_6604 <= p24_data_enable ? p23_bit_slice_6604 : p24_bit_slice_6604;
      p24_bit_slice_6605 <= p24_data_enable ? p23_bit_slice_6605 : p24_bit_slice_6605;
      p24_bit_slice_6606 <= p24_data_enable ? p23_bit_slice_6606 : p24_bit_slice_6606;
      p24_bit_slice_6607 <= p24_data_enable ? p23_bit_slice_6607 : p24_bit_slice_6607;
      p24_negated <= p24_data_enable ? p23_negated : p24_negated;
      p25_b <= p25_data_enable ? p24_b : p25_b;
      p25_uge_6683 <= p25_data_enable ? p24_uge_6683 : p25_uge_6683;
      p25_bivisor__1 <= p25_data_enable ? p24_bivisor__1 : p25_bivisor__1;
      p25_uge_6691 <= p25_data_enable ? p24_uge_6691 : p25_uge_6691;
      p25_uge_6771 <= p25_data_enable ? p24_uge_6771 : p25_uge_6771;
      p25_uge_6851 <= p25_data_enable ? p24_uge_6851 : p25_uge_6851;
      p25_uge_6931 <= p25_data_enable ? p24_uge_6931 : p25_uge_6931;
      p25_uge_7011 <= p25_data_enable ? p24_uge_7011 : p25_uge_7011;
      p25_uge_7091 <= p25_data_enable ? p24_uge_7091 : p25_uge_7091;
      p25_uge_7171 <= p25_data_enable ? p24_uge_7171 : p25_uge_7171;
      p25_uge_7251 <= p25_data_enable ? p24_uge_7251 : p25_uge_7251;
      p25_uge_7331 <= p25_data_enable ? p24_uge_7331 : p25_uge_7331;
      p25_uge_7411 <= p25_data_enable ? p24_uge_7411 : p25_uge_7411;
      p25_uge_7491 <= p25_data_enable ? p24_uge_7491 : p25_uge_7491;
      p25_uge_7571 <= p25_data_enable ? p24_uge_7571 : p25_uge_7571;
      p25_uge_7651 <= p25_data_enable ? p24_uge_7651 : p25_uge_7651;
      p25_uge_7731 <= p25_data_enable ? p24_uge_7731 : p25_uge_7731;
      p25_uge_7811 <= p25_data_enable ? p24_uge_7811 : p25_uge_7811;
      p25_uge_7891 <= p25_data_enable ? p24_uge_7891 : p25_uge_7891;
      p25_uge_7971 <= p25_data_enable ? p24_uge_7971 : p25_uge_7971;
      p25_uge_8051 <= p25_data_enable ? p24_uge_8051 : p25_uge_8051;
      p25_uge_8131 <= p25_data_enable ? p24_uge_8131 : p25_uge_8131;
      p25_uge_8211 <= p25_data_enable ? p24_uge_8211 : p25_uge_8211;
      p25_uge_8291 <= p25_data_enable ? p24_uge_8291 : p25_uge_8291;
      p25_uge_8371 <= p25_data_enable ? p24_uge_8371 : p25_uge_8371;
      p25_uge_8451 <= p25_data_enable ? p24_uge_8451 : p25_uge_8451;
      p25_uge_8531 <= p25_data_enable ? p24_uge_8531 : p25_uge_8531;
      p25_concat_8610 <= p25_data_enable ? concat_8610 : p25_concat_8610;
      p25_uge_8611 <= p25_data_enable ? uge_8611 : p25_uge_8611;
      p25_bit_slice_6602 <= p25_data_enable ? p24_bit_slice_6602 : p25_bit_slice_6602;
      p25_bit_slice_6603 <= p25_data_enable ? p24_bit_slice_6603 : p25_bit_slice_6603;
      p25_bit_slice_6604 <= p25_data_enable ? p24_bit_slice_6604 : p25_bit_slice_6604;
      p25_bit_slice_6605 <= p25_data_enable ? p24_bit_slice_6605 : p25_bit_slice_6605;
      p25_bit_slice_6606 <= p25_data_enable ? p24_bit_slice_6606 : p25_bit_slice_6606;
      p25_bit_slice_6607 <= p25_data_enable ? p24_bit_slice_6607 : p25_bit_slice_6607;
      p25_negated <= p25_data_enable ? p24_negated : p25_negated;
      p26_b <= p26_data_enable ? p25_b : p26_b;
      p26_uge_6683 <= p26_data_enable ? p25_uge_6683 : p26_uge_6683;
      p26_bivisor__1 <= p26_data_enable ? p25_bivisor__1 : p26_bivisor__1;
      p26_uge_6691 <= p26_data_enable ? p25_uge_6691 : p26_uge_6691;
      p26_uge_6771 <= p26_data_enable ? p25_uge_6771 : p26_uge_6771;
      p26_uge_6851 <= p26_data_enable ? p25_uge_6851 : p26_uge_6851;
      p26_uge_6931 <= p26_data_enable ? p25_uge_6931 : p26_uge_6931;
      p26_uge_7011 <= p26_data_enable ? p25_uge_7011 : p26_uge_7011;
      p26_uge_7091 <= p26_data_enable ? p25_uge_7091 : p26_uge_7091;
      p26_uge_7171 <= p26_data_enable ? p25_uge_7171 : p26_uge_7171;
      p26_uge_7251 <= p26_data_enable ? p25_uge_7251 : p26_uge_7251;
      p26_uge_7331 <= p26_data_enable ? p25_uge_7331 : p26_uge_7331;
      p26_uge_7411 <= p26_data_enable ? p25_uge_7411 : p26_uge_7411;
      p26_uge_7491 <= p26_data_enable ? p25_uge_7491 : p26_uge_7491;
      p26_uge_7571 <= p26_data_enable ? p25_uge_7571 : p26_uge_7571;
      p26_uge_7651 <= p26_data_enable ? p25_uge_7651 : p26_uge_7651;
      p26_uge_7731 <= p26_data_enable ? p25_uge_7731 : p26_uge_7731;
      p26_uge_7811 <= p26_data_enable ? p25_uge_7811 : p26_uge_7811;
      p26_uge_7891 <= p26_data_enable ? p25_uge_7891 : p26_uge_7891;
      p26_uge_7971 <= p26_data_enable ? p25_uge_7971 : p26_uge_7971;
      p26_uge_8051 <= p26_data_enable ? p25_uge_8051 : p26_uge_8051;
      p26_uge_8131 <= p26_data_enable ? p25_uge_8131 : p26_uge_8131;
      p26_uge_8211 <= p26_data_enable ? p25_uge_8211 : p26_uge_8211;
      p26_uge_8291 <= p26_data_enable ? p25_uge_8291 : p26_uge_8291;
      p26_uge_8371 <= p26_data_enable ? p25_uge_8371 : p26_uge_8371;
      p26_uge_8451 <= p26_data_enable ? p25_uge_8451 : p26_uge_8451;
      p26_uge_8531 <= p26_data_enable ? p25_uge_8531 : p26_uge_8531;
      p26_uge_8611 <= p26_data_enable ? p25_uge_8611 : p26_uge_8611;
      p26_concat_8690 <= p26_data_enable ? concat_8690 : p26_concat_8690;
      p26_uge_8691 <= p26_data_enable ? uge_8691 : p26_uge_8691;
      p26_bit_slice_6603 <= p26_data_enable ? p25_bit_slice_6603 : p26_bit_slice_6603;
      p26_bit_slice_6604 <= p26_data_enable ? p25_bit_slice_6604 : p26_bit_slice_6604;
      p26_bit_slice_6605 <= p26_data_enable ? p25_bit_slice_6605 : p26_bit_slice_6605;
      p26_bit_slice_6606 <= p26_data_enable ? p25_bit_slice_6606 : p26_bit_slice_6606;
      p26_bit_slice_6607 <= p26_data_enable ? p25_bit_slice_6607 : p26_bit_slice_6607;
      p26_negated <= p26_data_enable ? p25_negated : p26_negated;
      p27_b <= p27_data_enable ? p26_b : p27_b;
      p27_uge_6683 <= p27_data_enable ? p26_uge_6683 : p27_uge_6683;
      p27_bivisor__1 <= p27_data_enable ? p26_bivisor__1 : p27_bivisor__1;
      p27_uge_6691 <= p27_data_enable ? p26_uge_6691 : p27_uge_6691;
      p27_uge_6771 <= p27_data_enable ? p26_uge_6771 : p27_uge_6771;
      p27_uge_6851 <= p27_data_enable ? p26_uge_6851 : p27_uge_6851;
      p27_uge_6931 <= p27_data_enable ? p26_uge_6931 : p27_uge_6931;
      p27_uge_7011 <= p27_data_enable ? p26_uge_7011 : p27_uge_7011;
      p27_uge_7091 <= p27_data_enable ? p26_uge_7091 : p27_uge_7091;
      p27_uge_7171 <= p27_data_enable ? p26_uge_7171 : p27_uge_7171;
      p27_uge_7251 <= p27_data_enable ? p26_uge_7251 : p27_uge_7251;
      p27_uge_7331 <= p27_data_enable ? p26_uge_7331 : p27_uge_7331;
      p27_uge_7411 <= p27_data_enable ? p26_uge_7411 : p27_uge_7411;
      p27_uge_7491 <= p27_data_enable ? p26_uge_7491 : p27_uge_7491;
      p27_uge_7571 <= p27_data_enable ? p26_uge_7571 : p27_uge_7571;
      p27_uge_7651 <= p27_data_enable ? p26_uge_7651 : p27_uge_7651;
      p27_uge_7731 <= p27_data_enable ? p26_uge_7731 : p27_uge_7731;
      p27_uge_7811 <= p27_data_enable ? p26_uge_7811 : p27_uge_7811;
      p27_uge_7891 <= p27_data_enable ? p26_uge_7891 : p27_uge_7891;
      p27_uge_7971 <= p27_data_enable ? p26_uge_7971 : p27_uge_7971;
      p27_uge_8051 <= p27_data_enable ? p26_uge_8051 : p27_uge_8051;
      p27_uge_8131 <= p27_data_enable ? p26_uge_8131 : p27_uge_8131;
      p27_uge_8211 <= p27_data_enable ? p26_uge_8211 : p27_uge_8211;
      p27_uge_8291 <= p27_data_enable ? p26_uge_8291 : p27_uge_8291;
      p27_uge_8371 <= p27_data_enable ? p26_uge_8371 : p27_uge_8371;
      p27_uge_8451 <= p27_data_enable ? p26_uge_8451 : p27_uge_8451;
      p27_uge_8531 <= p27_data_enable ? p26_uge_8531 : p27_uge_8531;
      p27_uge_8611 <= p27_data_enable ? p26_uge_8611 : p27_uge_8611;
      p27_uge_8691 <= p27_data_enable ? p26_uge_8691 : p27_uge_8691;
      p27_concat_8770 <= p27_data_enable ? concat_8770 : p27_concat_8770;
      p27_uge_8771 <= p27_data_enable ? uge_8771 : p27_uge_8771;
      p27_bit_slice_6604 <= p27_data_enable ? p26_bit_slice_6604 : p27_bit_slice_6604;
      p27_bit_slice_6605 <= p27_data_enable ? p26_bit_slice_6605 : p27_bit_slice_6605;
      p27_bit_slice_6606 <= p27_data_enable ? p26_bit_slice_6606 : p27_bit_slice_6606;
      p27_bit_slice_6607 <= p27_data_enable ? p26_bit_slice_6607 : p27_bit_slice_6607;
      p27_negated <= p27_data_enable ? p26_negated : p27_negated;
      p28_b <= p28_data_enable ? p27_b : p28_b;
      p28_uge_6683 <= p28_data_enable ? p27_uge_6683 : p28_uge_6683;
      p28_bivisor__1 <= p28_data_enable ? p27_bivisor__1 : p28_bivisor__1;
      p28_uge_6691 <= p28_data_enable ? p27_uge_6691 : p28_uge_6691;
      p28_uge_6771 <= p28_data_enable ? p27_uge_6771 : p28_uge_6771;
      p28_uge_6851 <= p28_data_enable ? p27_uge_6851 : p28_uge_6851;
      p28_uge_6931 <= p28_data_enable ? p27_uge_6931 : p28_uge_6931;
      p28_uge_7011 <= p28_data_enable ? p27_uge_7011 : p28_uge_7011;
      p28_uge_7091 <= p28_data_enable ? p27_uge_7091 : p28_uge_7091;
      p28_uge_7171 <= p28_data_enable ? p27_uge_7171 : p28_uge_7171;
      p28_uge_7251 <= p28_data_enable ? p27_uge_7251 : p28_uge_7251;
      p28_uge_7331 <= p28_data_enable ? p27_uge_7331 : p28_uge_7331;
      p28_uge_7411 <= p28_data_enable ? p27_uge_7411 : p28_uge_7411;
      p28_uge_7491 <= p28_data_enable ? p27_uge_7491 : p28_uge_7491;
      p28_uge_7571 <= p28_data_enable ? p27_uge_7571 : p28_uge_7571;
      p28_uge_7651 <= p28_data_enable ? p27_uge_7651 : p28_uge_7651;
      p28_uge_7731 <= p28_data_enable ? p27_uge_7731 : p28_uge_7731;
      p28_uge_7811 <= p28_data_enable ? p27_uge_7811 : p28_uge_7811;
      p28_uge_7891 <= p28_data_enable ? p27_uge_7891 : p28_uge_7891;
      p28_uge_7971 <= p28_data_enable ? p27_uge_7971 : p28_uge_7971;
      p28_uge_8051 <= p28_data_enable ? p27_uge_8051 : p28_uge_8051;
      p28_uge_8131 <= p28_data_enable ? p27_uge_8131 : p28_uge_8131;
      p28_uge_8211 <= p28_data_enable ? p27_uge_8211 : p28_uge_8211;
      p28_uge_8291 <= p28_data_enable ? p27_uge_8291 : p28_uge_8291;
      p28_uge_8371 <= p28_data_enable ? p27_uge_8371 : p28_uge_8371;
      p28_uge_8451 <= p28_data_enable ? p27_uge_8451 : p28_uge_8451;
      p28_uge_8531 <= p28_data_enable ? p27_uge_8531 : p28_uge_8531;
      p28_uge_8611 <= p28_data_enable ? p27_uge_8611 : p28_uge_8611;
      p28_uge_8691 <= p28_data_enable ? p27_uge_8691 : p28_uge_8691;
      p28_uge_8771 <= p28_data_enable ? p27_uge_8771 : p28_uge_8771;
      p28_concat_8850 <= p28_data_enable ? concat_8850 : p28_concat_8850;
      p28_uge_8851 <= p28_data_enable ? uge_8851 : p28_uge_8851;
      p28_bit_slice_6605 <= p28_data_enable ? p27_bit_slice_6605 : p28_bit_slice_6605;
      p28_bit_slice_6606 <= p28_data_enable ? p27_bit_slice_6606 : p28_bit_slice_6606;
      p28_bit_slice_6607 <= p28_data_enable ? p27_bit_slice_6607 : p28_bit_slice_6607;
      p28_negated <= p28_data_enable ? p27_negated : p28_negated;
      p29_b <= p29_data_enable ? p28_b : p29_b;
      p29_uge_6683 <= p29_data_enable ? p28_uge_6683 : p29_uge_6683;
      p29_bivisor__1 <= p29_data_enable ? p28_bivisor__1 : p29_bivisor__1;
      p29_uge_6691 <= p29_data_enable ? p28_uge_6691 : p29_uge_6691;
      p29_uge_6771 <= p29_data_enable ? p28_uge_6771 : p29_uge_6771;
      p29_uge_6851 <= p29_data_enable ? p28_uge_6851 : p29_uge_6851;
      p29_uge_6931 <= p29_data_enable ? p28_uge_6931 : p29_uge_6931;
      p29_uge_7011 <= p29_data_enable ? p28_uge_7011 : p29_uge_7011;
      p29_uge_7091 <= p29_data_enable ? p28_uge_7091 : p29_uge_7091;
      p29_uge_7171 <= p29_data_enable ? p28_uge_7171 : p29_uge_7171;
      p29_uge_7251 <= p29_data_enable ? p28_uge_7251 : p29_uge_7251;
      p29_uge_7331 <= p29_data_enable ? p28_uge_7331 : p29_uge_7331;
      p29_uge_7411 <= p29_data_enable ? p28_uge_7411 : p29_uge_7411;
      p29_uge_7491 <= p29_data_enable ? p28_uge_7491 : p29_uge_7491;
      p29_uge_7571 <= p29_data_enable ? p28_uge_7571 : p29_uge_7571;
      p29_uge_7651 <= p29_data_enable ? p28_uge_7651 : p29_uge_7651;
      p29_uge_7731 <= p29_data_enable ? p28_uge_7731 : p29_uge_7731;
      p29_uge_7811 <= p29_data_enable ? p28_uge_7811 : p29_uge_7811;
      p29_uge_7891 <= p29_data_enable ? p28_uge_7891 : p29_uge_7891;
      p29_uge_7971 <= p29_data_enable ? p28_uge_7971 : p29_uge_7971;
      p29_uge_8051 <= p29_data_enable ? p28_uge_8051 : p29_uge_8051;
      p29_uge_8131 <= p29_data_enable ? p28_uge_8131 : p29_uge_8131;
      p29_uge_8211 <= p29_data_enable ? p28_uge_8211 : p29_uge_8211;
      p29_uge_8291 <= p29_data_enable ? p28_uge_8291 : p29_uge_8291;
      p29_uge_8371 <= p29_data_enable ? p28_uge_8371 : p29_uge_8371;
      p29_uge_8451 <= p29_data_enable ? p28_uge_8451 : p29_uge_8451;
      p29_uge_8531 <= p29_data_enable ? p28_uge_8531 : p29_uge_8531;
      p29_uge_8611 <= p29_data_enable ? p28_uge_8611 : p29_uge_8611;
      p29_uge_8691 <= p29_data_enable ? p28_uge_8691 : p29_uge_8691;
      p29_uge_8771 <= p29_data_enable ? p28_uge_8771 : p29_uge_8771;
      p29_uge_8851 <= p29_data_enable ? p28_uge_8851 : p29_uge_8851;
      p29_concat_8930 <= p29_data_enable ? concat_8930 : p29_concat_8930;
      p29_uge_8931 <= p29_data_enable ? uge_8931 : p29_uge_8931;
      p29_bit_slice_6606 <= p29_data_enable ? p28_bit_slice_6606 : p29_bit_slice_6606;
      p29_bit_slice_6607 <= p29_data_enable ? p28_bit_slice_6607 : p29_bit_slice_6607;
      p29_negated <= p29_data_enable ? p28_negated : p29_negated;
      p30_b <= p30_data_enable ? p29_b : p30_b;
      p30_uge_6683 <= p30_data_enable ? p29_uge_6683 : p30_uge_6683;
      p30_bivisor__1 <= p30_data_enable ? p29_bivisor__1 : p30_bivisor__1;
      p30_uge_6691 <= p30_data_enable ? p29_uge_6691 : p30_uge_6691;
      p30_uge_6771 <= p30_data_enable ? p29_uge_6771 : p30_uge_6771;
      p30_uge_6851 <= p30_data_enable ? p29_uge_6851 : p30_uge_6851;
      p30_uge_6931 <= p30_data_enable ? p29_uge_6931 : p30_uge_6931;
      p30_uge_7011 <= p30_data_enable ? p29_uge_7011 : p30_uge_7011;
      p30_uge_7091 <= p30_data_enable ? p29_uge_7091 : p30_uge_7091;
      p30_uge_7171 <= p30_data_enable ? p29_uge_7171 : p30_uge_7171;
      p30_uge_7251 <= p30_data_enable ? p29_uge_7251 : p30_uge_7251;
      p30_uge_7331 <= p30_data_enable ? p29_uge_7331 : p30_uge_7331;
      p30_uge_7411 <= p30_data_enable ? p29_uge_7411 : p30_uge_7411;
      p30_uge_7491 <= p30_data_enable ? p29_uge_7491 : p30_uge_7491;
      p30_uge_7571 <= p30_data_enable ? p29_uge_7571 : p30_uge_7571;
      p30_uge_7651 <= p30_data_enable ? p29_uge_7651 : p30_uge_7651;
      p30_uge_7731 <= p30_data_enable ? p29_uge_7731 : p30_uge_7731;
      p30_uge_7811 <= p30_data_enable ? p29_uge_7811 : p30_uge_7811;
      p30_uge_7891 <= p30_data_enable ? p29_uge_7891 : p30_uge_7891;
      p30_uge_7971 <= p30_data_enable ? p29_uge_7971 : p30_uge_7971;
      p30_uge_8051 <= p30_data_enable ? p29_uge_8051 : p30_uge_8051;
      p30_uge_8131 <= p30_data_enable ? p29_uge_8131 : p30_uge_8131;
      p30_uge_8211 <= p30_data_enable ? p29_uge_8211 : p30_uge_8211;
      p30_uge_8291 <= p30_data_enable ? p29_uge_8291 : p30_uge_8291;
      p30_uge_8371 <= p30_data_enable ? p29_uge_8371 : p30_uge_8371;
      p30_uge_8451 <= p30_data_enable ? p29_uge_8451 : p30_uge_8451;
      p30_uge_8531 <= p30_data_enable ? p29_uge_8531 : p30_uge_8531;
      p30_uge_8611 <= p30_data_enable ? p29_uge_8611 : p30_uge_8611;
      p30_uge_8691 <= p30_data_enable ? p29_uge_8691 : p30_uge_8691;
      p30_uge_8771 <= p30_data_enable ? p29_uge_8771 : p30_uge_8771;
      p30_uge_8851 <= p30_data_enable ? p29_uge_8851 : p30_uge_8851;
      p30_uge_8931 <= p30_data_enable ? p29_uge_8931 : p30_uge_8931;
      p30_concat_9010 <= p30_data_enable ? concat_9010 : p30_concat_9010;
      p30_uge_9011 <= p30_data_enable ? uge_9011 : p30_uge_9011;
      p30_bit_slice_6607 <= p30_data_enable ? p29_bit_slice_6607 : p30_bit_slice_6607;
      p30_negated <= p30_data_enable ? p29_negated : p30_negated;
      p31_uge_6683 <= p31_data_enable ? p30_uge_6683 : p31_uge_6683;
      p31_uge_6691 <= p31_data_enable ? p30_uge_6691 : p31_uge_6691;
      p31_uge_6771 <= p31_data_enable ? p30_uge_6771 : p31_uge_6771;
      p31_uge_6851 <= p31_data_enable ? p30_uge_6851 : p31_uge_6851;
      p31_uge_6931 <= p31_data_enable ? p30_uge_6931 : p31_uge_6931;
      p31_uge_7011 <= p31_data_enable ? p30_uge_7011 : p31_uge_7011;
      p31_uge_7091 <= p31_data_enable ? p30_uge_7091 : p31_uge_7091;
      p31_uge_7171 <= p31_data_enable ? p30_uge_7171 : p31_uge_7171;
      p31_uge_7251 <= p31_data_enable ? p30_uge_7251 : p31_uge_7251;
      p31_uge_7331 <= p31_data_enable ? p30_uge_7331 : p31_uge_7331;
      p31_uge_7411 <= p31_data_enable ? p30_uge_7411 : p31_uge_7411;
      p31_uge_7491 <= p31_data_enable ? p30_uge_7491 : p31_uge_7491;
      p31_uge_7571 <= p31_data_enable ? p30_uge_7571 : p31_uge_7571;
      p31_uge_7651 <= p31_data_enable ? p30_uge_7651 : p31_uge_7651;
      p31_uge_7731 <= p31_data_enable ? p30_uge_7731 : p31_uge_7731;
      p31_uge_7811 <= p31_data_enable ? p30_uge_7811 : p31_uge_7811;
      p31_uge_7891 <= p31_data_enable ? p30_uge_7891 : p31_uge_7891;
      p31_uge_7971 <= p31_data_enable ? p30_uge_7971 : p31_uge_7971;
      p31_uge_8051 <= p31_data_enable ? p30_uge_8051 : p31_uge_8051;
      p31_uge_8131 <= p31_data_enable ? p30_uge_8131 : p31_uge_8131;
      p31_uge_8211 <= p31_data_enable ? p30_uge_8211 : p31_uge_8211;
      p31_uge_8291 <= p31_data_enable ? p30_uge_8291 : p31_uge_8291;
      p31_uge_8371 <= p31_data_enable ? p30_uge_8371 : p31_uge_8371;
      p31_uge_8451 <= p31_data_enable ? p30_uge_8451 : p31_uge_8451;
      p31_uge_8531 <= p31_data_enable ? p30_uge_8531 : p31_uge_8531;
      p31_uge_8611 <= p31_data_enable ? p30_uge_8611 : p31_uge_8611;
      p31_uge_8691 <= p31_data_enable ? p30_uge_8691 : p31_uge_8691;
      p31_uge_8771 <= p31_data_enable ? p30_uge_8771 : p31_uge_8771;
      p31_uge_8851 <= p31_data_enable ? p30_uge_8851 : p31_uge_8851;
      p31_uge_8931 <= p31_data_enable ? p30_uge_8931 : p31_uge_8931;
      p31_uge_9011 <= p31_data_enable ? p30_uge_9011 : p31_uge_9011;
      p31_q__32_squeezed_portion_0_width_1 <= p31_data_enable ? q__32_squeezed_portion_0_width_1 : p31_q__32_squeezed_portion_0_width_1;
      p31_negated <= p31_data_enable ? p30_negated : p31_negated;
      p0_valid <= p0_enable ? p0_all_active_inputs_valid : p0_valid;
      p1_valid <= p1_enable ? p0_valid : p1_valid;
      p2_valid <= p2_enable ? p1_valid : p2_valid;
      p3_valid <= p3_enable ? p2_valid : p3_valid;
      p4_valid <= p4_enable ? p3_valid : p4_valid;
      p5_valid <= p5_enable ? p4_valid : p5_valid;
      p6_valid <= p6_enable ? p5_valid : p6_valid;
      p7_valid <= p7_enable ? p6_valid : p7_valid;
      p8_valid <= p8_enable ? p7_valid : p8_valid;
      p9_valid <= p9_enable ? p8_valid : p9_valid;
      p10_valid <= p10_enable ? p9_valid : p10_valid;
      p11_valid <= p11_enable ? p10_valid : p11_valid;
      p12_valid <= p12_enable ? p11_valid : p12_valid;
      p13_valid <= p13_enable ? p12_valid : p13_valid;
      p14_valid <= p14_enable ? p13_valid : p14_valid;
      p15_valid <= p15_enable ? p14_valid : p15_valid;
      p16_valid <= p16_enable ? p15_valid : p16_valid;
      p17_valid <= p17_enable ? p16_valid : p17_valid;
      p18_valid <= p18_enable ? p17_valid : p18_valid;
      p19_valid <= p19_enable ? p18_valid : p19_valid;
      p20_valid <= p20_enable ? p19_valid : p20_valid;
      p21_valid <= p21_enable ? p20_valid : p21_valid;
      p22_valid <= p22_enable ? p21_valid : p22_valid;
      p23_valid <= p23_enable ? p22_valid : p23_valid;
      p24_valid <= p24_enable ? p23_valid : p24_valid;
      p25_valid <= p25_enable ? p24_valid : p25_valid;
      p26_valid <= p26_enable ? p25_valid : p26_valid;
      p27_valid <= p27_enable ? p26_valid : p27_valid;
      p28_valid <= p28_enable ? p27_valid : p28_valid;
      p29_valid <= p29_enable ? p28_valid : p29_valid;
      p30_valid <= p30_enable ? p29_valid : p30_valid;
      p31_valid <= p31_enable ? p30_valid : p31_valid;
      p32_valid <= p32_enable ? p32_stage_done : p32_valid;
      p33_valid <= p33_enable ? p32_valid : p33_valid;
      p34_valid <= p34_enable ? p33_valid : p34_valid;
      __xls_float_ips__result_reg <= xls_float_ips__result_load_en ? __xls_float_ips__result_buf : __xls_float_ips__result_reg;
      __xls_float_ips__result_valid_reg <= xls_float_ips__result_valid_load_en ? p31_valid : __xls_float_ips__result_valid_reg;
    end
  end
  assign xls_float_ips__result = __xls_float_ips__result_reg;
  assign xls_float_ips__result_vld = __xls_float_ips__result_valid_reg;
  assign xls_float_ips__lhs_rdy = p0_data_enable;
  assign xls_float_ips__rhs_rdy = p0_data_enable;
endmodule
module __xls_float_ips__divui32_0_next(
  input wire clk,
  input wire rst,
  input wire [31:0] xls_float_ips__lhs,
  input wire xls_float_ips__lhs_vld,
  input wire [31:0] xls_float_ips__rhs,
  input wire xls_float_ips__rhs_vld,
  input wire xls_float_ips__result_rdy,
  output wire [31:0] xls_float_ips__result,
  output wire xls_float_ips__result_vld,
  output wire xls_float_ips__lhs_rdy,
  output wire xls_float_ips__rhs_rdy
);
  reg p0_bit_slice_6544;
  reg p0_bit_slice_6545;
  reg p0_bit_slice_6546;
  reg p0_bit_slice_6547;
  reg p0_bit_slice_6548;
  reg p0_bit_slice_6549;
  reg p0_bit_slice_6550;
  reg p0_bit_slice_6551;
  reg p0_bit_slice_6552;
  reg p0_bit_slice_6553;
  reg p0_bit_slice_6554;
  reg p0_bit_slice_6555;
  reg p0_bit_slice_6556;
  reg p0_bit_slice_6557;
  reg p0_bit_slice_6558;
  reg p0_bit_slice_6559;
  reg p0_bit_slice_6560;
  reg p0_bit_slice_6561;
  reg p0_bit_slice_6562;
  reg p0_bit_slice_6563;
  reg p0_bit_slice_6564;
  reg p0_bit_slice_6565;
  reg p0_bit_slice_6566;
  reg p0_bit_slice_6567;
  reg p0_bit_slice_6568;
  reg p0_bit_slice_6569;
  reg p0_bit_slice_6570;
  reg p0_bit_slice_6571;
  reg p0_bit_slice_6572;
  reg p0_bit_slice_6573;
  reg p0_bit_slice_6574;
  reg p0_bit_slice_6575;
  reg [31:0] p1_b;
  reg p1_uge_6652;
  reg [31:0] p1_r__2;
  reg p1_bit_slice_6545;
  reg p1_bit_slice_6546;
  reg p1_bit_slice_6547;
  reg p1_bit_slice_6548;
  reg p1_bit_slice_6549;
  reg p1_bit_slice_6550;
  reg p1_bit_slice_6551;
  reg p1_bit_slice_6552;
  reg p1_bit_slice_6553;
  reg p1_bit_slice_6554;
  reg p1_bit_slice_6555;
  reg p1_bit_slice_6556;
  reg p1_bit_slice_6557;
  reg p1_bit_slice_6558;
  reg p1_bit_slice_6559;
  reg p1_bit_slice_6560;
  reg p1_bit_slice_6561;
  reg p1_bit_slice_6562;
  reg p1_bit_slice_6563;
  reg p1_bit_slice_6564;
  reg p1_bit_slice_6565;
  reg p1_bit_slice_6566;
  reg p1_bit_slice_6567;
  reg p1_bit_slice_6568;
  reg p1_bit_slice_6569;
  reg p1_bit_slice_6570;
  reg p1_bit_slice_6571;
  reg p1_bit_slice_6572;
  reg p1_bit_slice_6573;
  reg p1_bit_slice_6574;
  reg p1_bit_slice_6575;
  reg [31:0] p2_b;
  reg p2_uge_6652;
  reg [32:0] p2_bivisor__1;
  reg p2_uge_6732;
  reg [31:0] p2_r__4;
  reg p2_bit_slice_6546;
  reg p2_bit_slice_6547;
  reg p2_bit_slice_6548;
  reg p2_bit_slice_6549;
  reg p2_bit_slice_6550;
  reg p2_bit_slice_6551;
  reg p2_bit_slice_6552;
  reg p2_bit_slice_6553;
  reg p2_bit_slice_6554;
  reg p2_bit_slice_6555;
  reg p2_bit_slice_6556;
  reg p2_bit_slice_6557;
  reg p2_bit_slice_6558;
  reg p2_bit_slice_6559;
  reg p2_bit_slice_6560;
  reg p2_bit_slice_6561;
  reg p2_bit_slice_6562;
  reg p2_bit_slice_6563;
  reg p2_bit_slice_6564;
  reg p2_bit_slice_6565;
  reg p2_bit_slice_6566;
  reg p2_bit_slice_6567;
  reg p2_bit_slice_6568;
  reg p2_bit_slice_6569;
  reg p2_bit_slice_6570;
  reg p2_bit_slice_6571;
  reg p2_bit_slice_6572;
  reg p2_bit_slice_6573;
  reg p2_bit_slice_6574;
  reg p2_bit_slice_6575;
  reg [31:0] p3_b;
  reg p3_uge_6652;
  reg [32:0] p3_bivisor__1;
  reg p3_uge_6732;
  reg p3_uge_6810;
  reg [31:0] p3_r__6;
  reg p3_bit_slice_6547;
  reg p3_bit_slice_6548;
  reg p3_bit_slice_6549;
  reg p3_bit_slice_6550;
  reg p3_bit_slice_6551;
  reg p3_bit_slice_6552;
  reg p3_bit_slice_6553;
  reg p3_bit_slice_6554;
  reg p3_bit_slice_6555;
  reg p3_bit_slice_6556;
  reg p3_bit_slice_6557;
  reg p3_bit_slice_6558;
  reg p3_bit_slice_6559;
  reg p3_bit_slice_6560;
  reg p3_bit_slice_6561;
  reg p3_bit_slice_6562;
  reg p3_bit_slice_6563;
  reg p3_bit_slice_6564;
  reg p3_bit_slice_6565;
  reg p3_bit_slice_6566;
  reg p3_bit_slice_6567;
  reg p3_bit_slice_6568;
  reg p3_bit_slice_6569;
  reg p3_bit_slice_6570;
  reg p3_bit_slice_6571;
  reg p3_bit_slice_6572;
  reg p3_bit_slice_6573;
  reg p3_bit_slice_6574;
  reg p3_bit_slice_6575;
  reg [31:0] p4_b;
  reg p4_uge_6652;
  reg [32:0] p4_bivisor__1;
  reg p4_uge_6732;
  reg p4_uge_6810;
  reg p4_uge_6888;
  reg [31:0] p4_r__8;
  reg p4_bit_slice_6548;
  reg p4_bit_slice_6549;
  reg p4_bit_slice_6550;
  reg p4_bit_slice_6551;
  reg p4_bit_slice_6552;
  reg p4_bit_slice_6553;
  reg p4_bit_slice_6554;
  reg p4_bit_slice_6555;
  reg p4_bit_slice_6556;
  reg p4_bit_slice_6557;
  reg p4_bit_slice_6558;
  reg p4_bit_slice_6559;
  reg p4_bit_slice_6560;
  reg p4_bit_slice_6561;
  reg p4_bit_slice_6562;
  reg p4_bit_slice_6563;
  reg p4_bit_slice_6564;
  reg p4_bit_slice_6565;
  reg p4_bit_slice_6566;
  reg p4_bit_slice_6567;
  reg p4_bit_slice_6568;
  reg p4_bit_slice_6569;
  reg p4_bit_slice_6570;
  reg p4_bit_slice_6571;
  reg p4_bit_slice_6572;
  reg p4_bit_slice_6573;
  reg p4_bit_slice_6574;
  reg p4_bit_slice_6575;
  reg [31:0] p5_b;
  reg p5_uge_6652;
  reg [32:0] p5_bivisor__1;
  reg p5_uge_6732;
  reg p5_uge_6810;
  reg p5_uge_6888;
  reg p5_uge_6966;
  reg [31:0] p5_r__10;
  reg p5_bit_slice_6549;
  reg p5_bit_slice_6550;
  reg p5_bit_slice_6551;
  reg p5_bit_slice_6552;
  reg p5_bit_slice_6553;
  reg p5_bit_slice_6554;
  reg p5_bit_slice_6555;
  reg p5_bit_slice_6556;
  reg p5_bit_slice_6557;
  reg p5_bit_slice_6558;
  reg p5_bit_slice_6559;
  reg p5_bit_slice_6560;
  reg p5_bit_slice_6561;
  reg p5_bit_slice_6562;
  reg p5_bit_slice_6563;
  reg p5_bit_slice_6564;
  reg p5_bit_slice_6565;
  reg p5_bit_slice_6566;
  reg p5_bit_slice_6567;
  reg p5_bit_slice_6568;
  reg p5_bit_slice_6569;
  reg p5_bit_slice_6570;
  reg p5_bit_slice_6571;
  reg p5_bit_slice_6572;
  reg p5_bit_slice_6573;
  reg p5_bit_slice_6574;
  reg p5_bit_slice_6575;
  reg [31:0] p6_b;
  reg p6_uge_6652;
  reg [32:0] p6_bivisor__1;
  reg p6_uge_6732;
  reg p6_uge_6810;
  reg p6_uge_6888;
  reg p6_uge_6966;
  reg p6_uge_7044;
  reg [31:0] p6_r__12;
  reg p6_bit_slice_6550;
  reg p6_bit_slice_6551;
  reg p6_bit_slice_6552;
  reg p6_bit_slice_6553;
  reg p6_bit_slice_6554;
  reg p6_bit_slice_6555;
  reg p6_bit_slice_6556;
  reg p6_bit_slice_6557;
  reg p6_bit_slice_6558;
  reg p6_bit_slice_6559;
  reg p6_bit_slice_6560;
  reg p6_bit_slice_6561;
  reg p6_bit_slice_6562;
  reg p6_bit_slice_6563;
  reg p6_bit_slice_6564;
  reg p6_bit_slice_6565;
  reg p6_bit_slice_6566;
  reg p6_bit_slice_6567;
  reg p6_bit_slice_6568;
  reg p6_bit_slice_6569;
  reg p6_bit_slice_6570;
  reg p6_bit_slice_6571;
  reg p6_bit_slice_6572;
  reg p6_bit_slice_6573;
  reg p6_bit_slice_6574;
  reg p6_bit_slice_6575;
  reg [31:0] p7_b;
  reg p7_uge_6652;
  reg [32:0] p7_bivisor__1;
  reg p7_uge_6732;
  reg p7_uge_6810;
  reg p7_uge_6888;
  reg p7_uge_6966;
  reg p7_uge_7044;
  reg p7_uge_7122;
  reg [31:0] p7_r__14;
  reg p7_bit_slice_6551;
  reg p7_bit_slice_6552;
  reg p7_bit_slice_6553;
  reg p7_bit_slice_6554;
  reg p7_bit_slice_6555;
  reg p7_bit_slice_6556;
  reg p7_bit_slice_6557;
  reg p7_bit_slice_6558;
  reg p7_bit_slice_6559;
  reg p7_bit_slice_6560;
  reg p7_bit_slice_6561;
  reg p7_bit_slice_6562;
  reg p7_bit_slice_6563;
  reg p7_bit_slice_6564;
  reg p7_bit_slice_6565;
  reg p7_bit_slice_6566;
  reg p7_bit_slice_6567;
  reg p7_bit_slice_6568;
  reg p7_bit_slice_6569;
  reg p7_bit_slice_6570;
  reg p7_bit_slice_6571;
  reg p7_bit_slice_6572;
  reg p7_bit_slice_6573;
  reg p7_bit_slice_6574;
  reg p7_bit_slice_6575;
  reg [31:0] p8_b;
  reg p8_uge_6652;
  reg [32:0] p8_bivisor__1;
  reg p8_uge_6732;
  reg p8_uge_6810;
  reg p8_uge_6888;
  reg p8_uge_6966;
  reg p8_uge_7044;
  reg p8_uge_7122;
  reg p8_uge_7200;
  reg [31:0] p8_r__16;
  reg p8_bit_slice_6552;
  reg p8_bit_slice_6553;
  reg p8_bit_slice_6554;
  reg p8_bit_slice_6555;
  reg p8_bit_slice_6556;
  reg p8_bit_slice_6557;
  reg p8_bit_slice_6558;
  reg p8_bit_slice_6559;
  reg p8_bit_slice_6560;
  reg p8_bit_slice_6561;
  reg p8_bit_slice_6562;
  reg p8_bit_slice_6563;
  reg p8_bit_slice_6564;
  reg p8_bit_slice_6565;
  reg p8_bit_slice_6566;
  reg p8_bit_slice_6567;
  reg p8_bit_slice_6568;
  reg p8_bit_slice_6569;
  reg p8_bit_slice_6570;
  reg p8_bit_slice_6571;
  reg p8_bit_slice_6572;
  reg p8_bit_slice_6573;
  reg p8_bit_slice_6574;
  reg p8_bit_slice_6575;
  reg [31:0] p9_b;
  reg p9_uge_6652;
  reg [32:0] p9_bivisor__1;
  reg p9_uge_6732;
  reg p9_uge_6810;
  reg p9_uge_6888;
  reg p9_uge_6966;
  reg p9_uge_7044;
  reg p9_uge_7122;
  reg p9_uge_7200;
  reg p9_uge_7278;
  reg [31:0] p9_r__18;
  reg p9_bit_slice_6553;
  reg p9_bit_slice_6554;
  reg p9_bit_slice_6555;
  reg p9_bit_slice_6556;
  reg p9_bit_slice_6557;
  reg p9_bit_slice_6558;
  reg p9_bit_slice_6559;
  reg p9_bit_slice_6560;
  reg p9_bit_slice_6561;
  reg p9_bit_slice_6562;
  reg p9_bit_slice_6563;
  reg p9_bit_slice_6564;
  reg p9_bit_slice_6565;
  reg p9_bit_slice_6566;
  reg p9_bit_slice_6567;
  reg p9_bit_slice_6568;
  reg p9_bit_slice_6569;
  reg p9_bit_slice_6570;
  reg p9_bit_slice_6571;
  reg p9_bit_slice_6572;
  reg p9_bit_slice_6573;
  reg p9_bit_slice_6574;
  reg p9_bit_slice_6575;
  reg [31:0] p10_b;
  reg p10_uge_6652;
  reg [32:0] p10_bivisor__1;
  reg p10_uge_6732;
  reg p10_uge_6810;
  reg p10_uge_6888;
  reg p10_uge_6966;
  reg p10_uge_7044;
  reg p10_uge_7122;
  reg p10_uge_7200;
  reg p10_uge_7278;
  reg p10_uge_7356;
  reg [31:0] p10_r__20;
  reg p10_bit_slice_6554;
  reg p10_bit_slice_6555;
  reg p10_bit_slice_6556;
  reg p10_bit_slice_6557;
  reg p10_bit_slice_6558;
  reg p10_bit_slice_6559;
  reg p10_bit_slice_6560;
  reg p10_bit_slice_6561;
  reg p10_bit_slice_6562;
  reg p10_bit_slice_6563;
  reg p10_bit_slice_6564;
  reg p10_bit_slice_6565;
  reg p10_bit_slice_6566;
  reg p10_bit_slice_6567;
  reg p10_bit_slice_6568;
  reg p10_bit_slice_6569;
  reg p10_bit_slice_6570;
  reg p10_bit_slice_6571;
  reg p10_bit_slice_6572;
  reg p10_bit_slice_6573;
  reg p10_bit_slice_6574;
  reg p10_bit_slice_6575;
  reg [31:0] p11_b;
  reg p11_uge_6652;
  reg [32:0] p11_bivisor__1;
  reg p11_uge_6732;
  reg p11_uge_6810;
  reg p11_uge_6888;
  reg p11_uge_6966;
  reg p11_uge_7044;
  reg p11_uge_7122;
  reg p11_uge_7200;
  reg p11_uge_7278;
  reg p11_uge_7356;
  reg p11_uge_7434;
  reg [31:0] p11_r__22;
  reg p11_bit_slice_6555;
  reg p11_bit_slice_6556;
  reg p11_bit_slice_6557;
  reg p11_bit_slice_6558;
  reg p11_bit_slice_6559;
  reg p11_bit_slice_6560;
  reg p11_bit_slice_6561;
  reg p11_bit_slice_6562;
  reg p11_bit_slice_6563;
  reg p11_bit_slice_6564;
  reg p11_bit_slice_6565;
  reg p11_bit_slice_6566;
  reg p11_bit_slice_6567;
  reg p11_bit_slice_6568;
  reg p11_bit_slice_6569;
  reg p11_bit_slice_6570;
  reg p11_bit_slice_6571;
  reg p11_bit_slice_6572;
  reg p11_bit_slice_6573;
  reg p11_bit_slice_6574;
  reg p11_bit_slice_6575;
  reg [31:0] p12_b;
  reg p12_uge_6652;
  reg [32:0] p12_bivisor__1;
  reg p12_uge_6732;
  reg p12_uge_6810;
  reg p12_uge_6888;
  reg p12_uge_6966;
  reg p12_uge_7044;
  reg p12_uge_7122;
  reg p12_uge_7200;
  reg p12_uge_7278;
  reg p12_uge_7356;
  reg p12_uge_7434;
  reg p12_uge_7512;
  reg [31:0] p12_r__24;
  reg p12_bit_slice_6556;
  reg p12_bit_slice_6557;
  reg p12_bit_slice_6558;
  reg p12_bit_slice_6559;
  reg p12_bit_slice_6560;
  reg p12_bit_slice_6561;
  reg p12_bit_slice_6562;
  reg p12_bit_slice_6563;
  reg p12_bit_slice_6564;
  reg p12_bit_slice_6565;
  reg p12_bit_slice_6566;
  reg p12_bit_slice_6567;
  reg p12_bit_slice_6568;
  reg p12_bit_slice_6569;
  reg p12_bit_slice_6570;
  reg p12_bit_slice_6571;
  reg p12_bit_slice_6572;
  reg p12_bit_slice_6573;
  reg p12_bit_slice_6574;
  reg p12_bit_slice_6575;
  reg [31:0] p13_b;
  reg p13_uge_6652;
  reg [32:0] p13_bivisor__1;
  reg p13_uge_6732;
  reg p13_uge_6810;
  reg p13_uge_6888;
  reg p13_uge_6966;
  reg p13_uge_7044;
  reg p13_uge_7122;
  reg p13_uge_7200;
  reg p13_uge_7278;
  reg p13_uge_7356;
  reg p13_uge_7434;
  reg p13_uge_7512;
  reg p13_uge_7590;
  reg [31:0] p13_r__26;
  reg p13_bit_slice_6557;
  reg p13_bit_slice_6558;
  reg p13_bit_slice_6559;
  reg p13_bit_slice_6560;
  reg p13_bit_slice_6561;
  reg p13_bit_slice_6562;
  reg p13_bit_slice_6563;
  reg p13_bit_slice_6564;
  reg p13_bit_slice_6565;
  reg p13_bit_slice_6566;
  reg p13_bit_slice_6567;
  reg p13_bit_slice_6568;
  reg p13_bit_slice_6569;
  reg p13_bit_slice_6570;
  reg p13_bit_slice_6571;
  reg p13_bit_slice_6572;
  reg p13_bit_slice_6573;
  reg p13_bit_slice_6574;
  reg p13_bit_slice_6575;
  reg [31:0] p14_b;
  reg p14_uge_6652;
  reg [32:0] p14_bivisor__1;
  reg p14_uge_6732;
  reg p14_uge_6810;
  reg p14_uge_6888;
  reg p14_uge_6966;
  reg p14_uge_7044;
  reg p14_uge_7122;
  reg p14_uge_7200;
  reg p14_uge_7278;
  reg p14_uge_7356;
  reg p14_uge_7434;
  reg p14_uge_7512;
  reg p14_uge_7590;
  reg p14_uge_7668;
  reg [31:0] p14_r__28;
  reg p14_bit_slice_6558;
  reg p14_bit_slice_6559;
  reg p14_bit_slice_6560;
  reg p14_bit_slice_6561;
  reg p14_bit_slice_6562;
  reg p14_bit_slice_6563;
  reg p14_bit_slice_6564;
  reg p14_bit_slice_6565;
  reg p14_bit_slice_6566;
  reg p14_bit_slice_6567;
  reg p14_bit_slice_6568;
  reg p14_bit_slice_6569;
  reg p14_bit_slice_6570;
  reg p14_bit_slice_6571;
  reg p14_bit_slice_6572;
  reg p14_bit_slice_6573;
  reg p14_bit_slice_6574;
  reg p14_bit_slice_6575;
  reg [31:0] p15_b;
  reg p15_uge_6652;
  reg [32:0] p15_bivisor__1;
  reg p15_uge_6732;
  reg p15_uge_6810;
  reg p15_uge_6888;
  reg p15_uge_6966;
  reg p15_uge_7044;
  reg p15_uge_7122;
  reg p15_uge_7200;
  reg p15_uge_7278;
  reg p15_uge_7356;
  reg p15_uge_7434;
  reg p15_uge_7512;
  reg p15_uge_7590;
  reg p15_uge_7668;
  reg p15_uge_7746;
  reg [31:0] p15_r__30;
  reg p15_bit_slice_6559;
  reg p15_bit_slice_6560;
  reg p15_bit_slice_6561;
  reg p15_bit_slice_6562;
  reg p15_bit_slice_6563;
  reg p15_bit_slice_6564;
  reg p15_bit_slice_6565;
  reg p15_bit_slice_6566;
  reg p15_bit_slice_6567;
  reg p15_bit_slice_6568;
  reg p15_bit_slice_6569;
  reg p15_bit_slice_6570;
  reg p15_bit_slice_6571;
  reg p15_bit_slice_6572;
  reg p15_bit_slice_6573;
  reg p15_bit_slice_6574;
  reg p15_bit_slice_6575;
  reg [31:0] p16_b;
  reg p16_uge_6652;
  reg [32:0] p16_bivisor__1;
  reg p16_uge_6732;
  reg p16_uge_6810;
  reg p16_uge_6888;
  reg p16_uge_6966;
  reg p16_uge_7044;
  reg p16_uge_7122;
  reg p16_uge_7200;
  reg p16_uge_7278;
  reg p16_uge_7356;
  reg p16_uge_7434;
  reg p16_uge_7512;
  reg p16_uge_7590;
  reg p16_uge_7668;
  reg p16_uge_7746;
  reg p16_uge_7824;
  reg [31:0] p16_r__32;
  reg p16_bit_slice_6560;
  reg p16_bit_slice_6561;
  reg p16_bit_slice_6562;
  reg p16_bit_slice_6563;
  reg p16_bit_slice_6564;
  reg p16_bit_slice_6565;
  reg p16_bit_slice_6566;
  reg p16_bit_slice_6567;
  reg p16_bit_slice_6568;
  reg p16_bit_slice_6569;
  reg p16_bit_slice_6570;
  reg p16_bit_slice_6571;
  reg p16_bit_slice_6572;
  reg p16_bit_slice_6573;
  reg p16_bit_slice_6574;
  reg p16_bit_slice_6575;
  reg [31:0] p17_b;
  reg p17_uge_6652;
  reg [32:0] p17_bivisor__1;
  reg p17_uge_6732;
  reg p17_uge_6810;
  reg p17_uge_6888;
  reg p17_uge_6966;
  reg p17_uge_7044;
  reg p17_uge_7122;
  reg p17_uge_7200;
  reg p17_uge_7278;
  reg p17_uge_7356;
  reg p17_uge_7434;
  reg p17_uge_7512;
  reg p17_uge_7590;
  reg p17_uge_7668;
  reg p17_uge_7746;
  reg p17_uge_7824;
  reg p17_uge_7902;
  reg [31:0] p17_r__34;
  reg p17_bit_slice_6561;
  reg p17_bit_slice_6562;
  reg p17_bit_slice_6563;
  reg p17_bit_slice_6564;
  reg p17_bit_slice_6565;
  reg p17_bit_slice_6566;
  reg p17_bit_slice_6567;
  reg p17_bit_slice_6568;
  reg p17_bit_slice_6569;
  reg p17_bit_slice_6570;
  reg p17_bit_slice_6571;
  reg p17_bit_slice_6572;
  reg p17_bit_slice_6573;
  reg p17_bit_slice_6574;
  reg p17_bit_slice_6575;
  reg [31:0] p18_b;
  reg p18_uge_6652;
  reg [32:0] p18_bivisor__1;
  reg p18_uge_6732;
  reg p18_uge_6810;
  reg p18_uge_6888;
  reg p18_uge_6966;
  reg p18_uge_7044;
  reg p18_uge_7122;
  reg p18_uge_7200;
  reg p18_uge_7278;
  reg p18_uge_7356;
  reg p18_uge_7434;
  reg p18_uge_7512;
  reg p18_uge_7590;
  reg p18_uge_7668;
  reg p18_uge_7746;
  reg p18_uge_7824;
  reg p18_uge_7902;
  reg p18_uge_7980;
  reg [31:0] p18_r__36;
  reg p18_bit_slice_6562;
  reg p18_bit_slice_6563;
  reg p18_bit_slice_6564;
  reg p18_bit_slice_6565;
  reg p18_bit_slice_6566;
  reg p18_bit_slice_6567;
  reg p18_bit_slice_6568;
  reg p18_bit_slice_6569;
  reg p18_bit_slice_6570;
  reg p18_bit_slice_6571;
  reg p18_bit_slice_6572;
  reg p18_bit_slice_6573;
  reg p18_bit_slice_6574;
  reg p18_bit_slice_6575;
  reg [31:0] p19_b;
  reg p19_uge_6652;
  reg [32:0] p19_bivisor__1;
  reg p19_uge_6732;
  reg p19_uge_6810;
  reg p19_uge_6888;
  reg p19_uge_6966;
  reg p19_uge_7044;
  reg p19_uge_7122;
  reg p19_uge_7200;
  reg p19_uge_7278;
  reg p19_uge_7356;
  reg p19_uge_7434;
  reg p19_uge_7512;
  reg p19_uge_7590;
  reg p19_uge_7668;
  reg p19_uge_7746;
  reg p19_uge_7824;
  reg p19_uge_7902;
  reg p19_uge_7980;
  reg p19_uge_8058;
  reg [31:0] p19_r__38;
  reg p19_bit_slice_6563;
  reg p19_bit_slice_6564;
  reg p19_bit_slice_6565;
  reg p19_bit_slice_6566;
  reg p19_bit_slice_6567;
  reg p19_bit_slice_6568;
  reg p19_bit_slice_6569;
  reg p19_bit_slice_6570;
  reg p19_bit_slice_6571;
  reg p19_bit_slice_6572;
  reg p19_bit_slice_6573;
  reg p19_bit_slice_6574;
  reg p19_bit_slice_6575;
  reg [31:0] p20_b;
  reg p20_uge_6652;
  reg [32:0] p20_bivisor__1;
  reg p20_uge_6732;
  reg p20_uge_6810;
  reg p20_uge_6888;
  reg p20_uge_6966;
  reg p20_uge_7044;
  reg p20_uge_7122;
  reg p20_uge_7200;
  reg p20_uge_7278;
  reg p20_uge_7356;
  reg p20_uge_7434;
  reg p20_uge_7512;
  reg p20_uge_7590;
  reg p20_uge_7668;
  reg p20_uge_7746;
  reg p20_uge_7824;
  reg p20_uge_7902;
  reg p20_uge_7980;
  reg p20_uge_8058;
  reg p20_uge_8136;
  reg [31:0] p20_r__40;
  reg p20_bit_slice_6564;
  reg p20_bit_slice_6565;
  reg p20_bit_slice_6566;
  reg p20_bit_slice_6567;
  reg p20_bit_slice_6568;
  reg p20_bit_slice_6569;
  reg p20_bit_slice_6570;
  reg p20_bit_slice_6571;
  reg p20_bit_slice_6572;
  reg p20_bit_slice_6573;
  reg p20_bit_slice_6574;
  reg p20_bit_slice_6575;
  reg [31:0] p21_b;
  reg p21_uge_6652;
  reg [32:0] p21_bivisor__1;
  reg p21_uge_6732;
  reg p21_uge_6810;
  reg p21_uge_6888;
  reg p21_uge_6966;
  reg p21_uge_7044;
  reg p21_uge_7122;
  reg p21_uge_7200;
  reg p21_uge_7278;
  reg p21_uge_7356;
  reg p21_uge_7434;
  reg p21_uge_7512;
  reg p21_uge_7590;
  reg p21_uge_7668;
  reg p21_uge_7746;
  reg p21_uge_7824;
  reg p21_uge_7902;
  reg p21_uge_7980;
  reg p21_uge_8058;
  reg p21_uge_8136;
  reg p21_uge_8214;
  reg [31:0] p21_r__42;
  reg p21_bit_slice_6565;
  reg p21_bit_slice_6566;
  reg p21_bit_slice_6567;
  reg p21_bit_slice_6568;
  reg p21_bit_slice_6569;
  reg p21_bit_slice_6570;
  reg p21_bit_slice_6571;
  reg p21_bit_slice_6572;
  reg p21_bit_slice_6573;
  reg p21_bit_slice_6574;
  reg p21_bit_slice_6575;
  reg [31:0] p22_b;
  reg p22_uge_6652;
  reg [32:0] p22_bivisor__1;
  reg p22_uge_6732;
  reg p22_uge_6810;
  reg p22_uge_6888;
  reg p22_uge_6966;
  reg p22_uge_7044;
  reg p22_uge_7122;
  reg p22_uge_7200;
  reg p22_uge_7278;
  reg p22_uge_7356;
  reg p22_uge_7434;
  reg p22_uge_7512;
  reg p22_uge_7590;
  reg p22_uge_7668;
  reg p22_uge_7746;
  reg p22_uge_7824;
  reg p22_uge_7902;
  reg p22_uge_7980;
  reg p22_uge_8058;
  reg p22_uge_8136;
  reg p22_uge_8214;
  reg p22_uge_8292;
  reg [31:0] p22_r__44;
  reg p22_bit_slice_6566;
  reg p22_bit_slice_6567;
  reg p22_bit_slice_6568;
  reg p22_bit_slice_6569;
  reg p22_bit_slice_6570;
  reg p22_bit_slice_6571;
  reg p22_bit_slice_6572;
  reg p22_bit_slice_6573;
  reg p22_bit_slice_6574;
  reg p22_bit_slice_6575;
  reg [31:0] p23_b;
  reg p23_uge_6652;
  reg [32:0] p23_bivisor__1;
  reg p23_uge_6732;
  reg p23_uge_6810;
  reg p23_uge_6888;
  reg p23_uge_6966;
  reg p23_uge_7044;
  reg p23_uge_7122;
  reg p23_uge_7200;
  reg p23_uge_7278;
  reg p23_uge_7356;
  reg p23_uge_7434;
  reg p23_uge_7512;
  reg p23_uge_7590;
  reg p23_uge_7668;
  reg p23_uge_7746;
  reg p23_uge_7824;
  reg p23_uge_7902;
  reg p23_uge_7980;
  reg p23_uge_8058;
  reg p23_uge_8136;
  reg p23_uge_8214;
  reg p23_uge_8292;
  reg p23_uge_8370;
  reg [31:0] p23_r__46;
  reg p23_bit_slice_6567;
  reg p23_bit_slice_6568;
  reg p23_bit_slice_6569;
  reg p23_bit_slice_6570;
  reg p23_bit_slice_6571;
  reg p23_bit_slice_6572;
  reg p23_bit_slice_6573;
  reg p23_bit_slice_6574;
  reg p23_bit_slice_6575;
  reg [31:0] p24_b;
  reg p24_uge_6652;
  reg [32:0] p24_bivisor__1;
  reg p24_uge_6732;
  reg p24_uge_6810;
  reg p24_uge_6888;
  reg p24_uge_6966;
  reg p24_uge_7044;
  reg p24_uge_7122;
  reg p24_uge_7200;
  reg p24_uge_7278;
  reg p24_uge_7356;
  reg p24_uge_7434;
  reg p24_uge_7512;
  reg p24_uge_7590;
  reg p24_uge_7668;
  reg p24_uge_7746;
  reg p24_uge_7824;
  reg p24_uge_7902;
  reg p24_uge_7980;
  reg p24_uge_8058;
  reg p24_uge_8136;
  reg p24_uge_8214;
  reg p24_uge_8292;
  reg p24_uge_8370;
  reg p24_uge_8448;
  reg [31:0] p24_r__48;
  reg p24_bit_slice_6568;
  reg p24_bit_slice_6569;
  reg p24_bit_slice_6570;
  reg p24_bit_slice_6571;
  reg p24_bit_slice_6572;
  reg p24_bit_slice_6573;
  reg p24_bit_slice_6574;
  reg p24_bit_slice_6575;
  reg [31:0] p25_b;
  reg p25_uge_6652;
  reg [32:0] p25_bivisor__1;
  reg p25_uge_6732;
  reg p25_uge_6810;
  reg p25_uge_6888;
  reg p25_uge_6966;
  reg p25_uge_7044;
  reg p25_uge_7122;
  reg p25_uge_7200;
  reg p25_uge_7278;
  reg p25_uge_7356;
  reg p25_uge_7434;
  reg p25_uge_7512;
  reg p25_uge_7590;
  reg p25_uge_7668;
  reg p25_uge_7746;
  reg p25_uge_7824;
  reg p25_uge_7902;
  reg p25_uge_7980;
  reg p25_uge_8058;
  reg p25_uge_8136;
  reg p25_uge_8214;
  reg p25_uge_8292;
  reg p25_uge_8370;
  reg p25_uge_8448;
  reg p25_uge_8526;
  reg [31:0] p25_r__50;
  reg p25_bit_slice_6569;
  reg p25_bit_slice_6570;
  reg p25_bit_slice_6571;
  reg p25_bit_slice_6572;
  reg p25_bit_slice_6573;
  reg p25_bit_slice_6574;
  reg p25_bit_slice_6575;
  reg [31:0] p26_b;
  reg p26_uge_6652;
  reg [32:0] p26_bivisor__1;
  reg p26_uge_6732;
  reg p26_uge_6810;
  reg p26_uge_6888;
  reg p26_uge_6966;
  reg p26_uge_7044;
  reg p26_uge_7122;
  reg p26_uge_7200;
  reg p26_uge_7278;
  reg p26_uge_7356;
  reg p26_uge_7434;
  reg p26_uge_7512;
  reg p26_uge_7590;
  reg p26_uge_7668;
  reg p26_uge_7746;
  reg p26_uge_7824;
  reg p26_uge_7902;
  reg p26_uge_7980;
  reg p26_uge_8058;
  reg p26_uge_8136;
  reg p26_uge_8214;
  reg p26_uge_8292;
  reg p26_uge_8370;
  reg p26_uge_8448;
  reg p26_uge_8526;
  reg p26_uge_8604;
  reg [31:0] p26_r__52;
  reg p26_bit_slice_6570;
  reg p26_bit_slice_6571;
  reg p26_bit_slice_6572;
  reg p26_bit_slice_6573;
  reg p26_bit_slice_6574;
  reg p26_bit_slice_6575;
  reg [31:0] p27_b;
  reg p27_uge_6652;
  reg [32:0] p27_bivisor__1;
  reg p27_uge_6732;
  reg p27_uge_6810;
  reg p27_uge_6888;
  reg p27_uge_6966;
  reg p27_uge_7044;
  reg p27_uge_7122;
  reg p27_uge_7200;
  reg p27_uge_7278;
  reg p27_uge_7356;
  reg p27_uge_7434;
  reg p27_uge_7512;
  reg p27_uge_7590;
  reg p27_uge_7668;
  reg p27_uge_7746;
  reg p27_uge_7824;
  reg p27_uge_7902;
  reg p27_uge_7980;
  reg p27_uge_8058;
  reg p27_uge_8136;
  reg p27_uge_8214;
  reg p27_uge_8292;
  reg p27_uge_8370;
  reg p27_uge_8448;
  reg p27_uge_8526;
  reg p27_uge_8604;
  reg p27_uge_8682;
  reg [31:0] p27_r__54;
  reg p27_bit_slice_6571;
  reg p27_bit_slice_6572;
  reg p27_bit_slice_6573;
  reg p27_bit_slice_6574;
  reg p27_bit_slice_6575;
  reg [31:0] p28_b;
  reg p28_uge_6652;
  reg [32:0] p28_bivisor__1;
  reg p28_uge_6732;
  reg p28_uge_6810;
  reg p28_uge_6888;
  reg p28_uge_6966;
  reg p28_uge_7044;
  reg p28_uge_7122;
  reg p28_uge_7200;
  reg p28_uge_7278;
  reg p28_uge_7356;
  reg p28_uge_7434;
  reg p28_uge_7512;
  reg p28_uge_7590;
  reg p28_uge_7668;
  reg p28_uge_7746;
  reg p28_uge_7824;
  reg p28_uge_7902;
  reg p28_uge_7980;
  reg p28_uge_8058;
  reg p28_uge_8136;
  reg p28_uge_8214;
  reg p28_uge_8292;
  reg p28_uge_8370;
  reg p28_uge_8448;
  reg p28_uge_8526;
  reg p28_uge_8604;
  reg p28_uge_8682;
  reg p28_uge_8760;
  reg [31:0] p28_r__56;
  reg p28_bit_slice_6572;
  reg p28_bit_slice_6573;
  reg p28_bit_slice_6574;
  reg p28_bit_slice_6575;
  reg [31:0] p29_b;
  reg p29_uge_6652;
  reg [32:0] p29_bivisor__1;
  reg p29_uge_6732;
  reg p29_uge_6810;
  reg p29_uge_6888;
  reg p29_uge_6966;
  reg p29_uge_7044;
  reg p29_uge_7122;
  reg p29_uge_7200;
  reg p29_uge_7278;
  reg p29_uge_7356;
  reg p29_uge_7434;
  reg p29_uge_7512;
  reg p29_uge_7590;
  reg p29_uge_7668;
  reg p29_uge_7746;
  reg p29_uge_7824;
  reg p29_uge_7902;
  reg p29_uge_7980;
  reg p29_uge_8058;
  reg p29_uge_8136;
  reg p29_uge_8214;
  reg p29_uge_8292;
  reg p29_uge_8370;
  reg p29_uge_8448;
  reg p29_uge_8526;
  reg p29_uge_8604;
  reg p29_uge_8682;
  reg p29_uge_8760;
  reg p29_uge_8838;
  reg [31:0] p29_r__58;
  reg p29_bit_slice_6573;
  reg p29_bit_slice_6574;
  reg p29_bit_slice_6575;
  reg [31:0] p30_b;
  reg p30_uge_6652;
  reg [32:0] p30_bivisor__1;
  reg p30_uge_6732;
  reg p30_uge_6810;
  reg p30_uge_6888;
  reg p30_uge_6966;
  reg p30_uge_7044;
  reg p30_uge_7122;
  reg p30_uge_7200;
  reg p30_uge_7278;
  reg p30_uge_7356;
  reg p30_uge_7434;
  reg p30_uge_7512;
  reg p30_uge_7590;
  reg p30_uge_7668;
  reg p30_uge_7746;
  reg p30_uge_7824;
  reg p30_uge_7902;
  reg p30_uge_7980;
  reg p30_uge_8058;
  reg p30_uge_8136;
  reg p30_uge_8214;
  reg p30_uge_8292;
  reg p30_uge_8370;
  reg p30_uge_8448;
  reg p30_uge_8526;
  reg p30_uge_8604;
  reg p30_uge_8682;
  reg p30_uge_8760;
  reg p30_uge_8838;
  reg p30_uge_8916;
  reg [31:0] p30_r__60;
  reg p30_bit_slice_6574;
  reg p30_bit_slice_6575;
  reg p31_uge_6652;
  reg [32:0] p31_bivisor__1;
  reg p31_uge_6732;
  reg p31_uge_6810;
  reg p31_uge_6888;
  reg p31_uge_6966;
  reg p31_uge_7044;
  reg p31_uge_7122;
  reg p31_uge_7200;
  reg p31_uge_7278;
  reg p31_uge_7356;
  reg p31_uge_7434;
  reg p31_uge_7512;
  reg p31_uge_7590;
  reg p31_uge_7668;
  reg p31_uge_7746;
  reg p31_uge_7824;
  reg p31_uge_7902;
  reg p31_uge_7980;
  reg p31_uge_8058;
  reg p31_uge_8136;
  reg p31_uge_8214;
  reg p31_uge_8292;
  reg p31_uge_8370;
  reg p31_uge_8448;
  reg p31_uge_8526;
  reg p31_uge_8604;
  reg p31_uge_8682;
  reg p31_uge_8760;
  reg p31_uge_8838;
  reg p31_uge_8916;
  reg p31_uge_8994;
  reg [31:0] p31_r__62;
  reg p31_bit_slice_6575;
  reg p0_valid;
  reg p1_valid;
  reg p2_valid;
  reg p3_valid;
  reg p4_valid;
  reg p5_valid;
  reg p6_valid;
  reg p7_valid;
  reg p8_valid;
  reg p9_valid;
  reg p10_valid;
  reg p11_valid;
  reg p12_valid;
  reg p13_valid;
  reg p14_valid;
  reg p15_valid;
  reg p16_valid;
  reg p17_valid;
  reg p18_valid;
  reg p19_valid;
  reg p20_valid;
  reg p21_valid;
  reg p22_valid;
  reg p23_valid;
  reg p24_valid;
  reg p25_valid;
  reg p26_valid;
  reg p27_valid;
  reg p28_valid;
  reg p29_valid;
  reg p30_valid;
  reg p31_valid;
  reg p32_valid;
  reg p33_valid;
  reg p34_valid;
  reg [31:0] __xls_float_ips__result_reg;
  reg __xls_float_ips__result_valid_reg;
  wire xls_float_ips__result_valid_inv;
  wire xls_float_ips__result_valid_load_en;
  wire xls_float_ips__result_load_en;
  wire p32_stage_done;
  wire p32_not_valid;
  wire p31_enable;
  wire p31_data_enable;
  wire p31_not_valid;
  wire p30_enable;
  wire p30_data_enable;
  wire p30_not_valid;
  wire p29_enable;
  wire p29_data_enable;
  wire p29_not_valid;
  wire p28_enable;
  wire p28_data_enable;
  wire p28_not_valid;
  wire p27_enable;
  wire p27_data_enable;
  wire p27_not_valid;
  wire p26_enable;
  wire p26_data_enable;
  wire p26_not_valid;
  wire p25_enable;
  wire p25_data_enable;
  wire p25_not_valid;
  wire p24_enable;
  wire p24_data_enable;
  wire p24_not_valid;
  wire p23_enable;
  wire p23_data_enable;
  wire p23_not_valid;
  wire p22_enable;
  wire p22_data_enable;
  wire p22_not_valid;
  wire p21_enable;
  wire p21_data_enable;
  wire p21_not_valid;
  wire p20_enable;
  wire p20_data_enable;
  wire p20_not_valid;
  wire p19_enable;
  wire p19_data_enable;
  wire p19_not_valid;
  wire p18_enable;
  wire p18_data_enable;
  wire p18_not_valid;
  wire p17_enable;
  wire p17_data_enable;
  wire p17_not_valid;
  wire p16_enable;
  wire p16_data_enable;
  wire p16_not_valid;
  wire p15_enable;
  wire p15_data_enable;
  wire p15_not_valid;
  wire p14_enable;
  wire p14_data_enable;
  wire p14_not_valid;
  wire p13_enable;
  wire p13_data_enable;
  wire p13_not_valid;
  wire p12_enable;
  wire p12_data_enable;
  wire p12_not_valid;
  wire p11_enable;
  wire p11_data_enable;
  wire p11_not_valid;
  wire p10_enable;
  wire p10_data_enable;
  wire p10_not_valid;
  wire p9_enable;
  wire p9_data_enable;
  wire p9_not_valid;
  wire p8_enable;
  wire p8_data_enable;
  wire p8_not_valid;
  wire p7_enable;
  wire p7_data_enable;
  wire p7_not_valid;
  wire p6_enable;
  wire p6_data_enable;
  wire p6_not_valid;
  wire p5_enable;
  wire p5_data_enable;
  wire p5_not_valid;
  wire p4_enable;
  wire p4_data_enable;
  wire p4_not_valid;
  wire p3_enable;
  wire p3_data_enable;
  wire p3_not_valid;
  wire p2_enable;
  wire p2_data_enable;
  wire p2_not_valid;
  wire p1_enable;
  wire p1_stage_done;
  wire [32:0] r__61;
  wire [31:0] concat_8993;
  wire [32:0] r__59;
  wire [31:0] concat_8915;
  wire [32:0] r__57;
  wire [31:0] concat_8837;
  wire [32:0] r__55;
  wire [31:0] concat_8759;
  wire [32:0] r__53;
  wire [31:0] concat_8681;
  wire [32:0] r__51;
  wire [31:0] concat_8603;
  wire [32:0] r__49;
  wire [31:0] concat_8525;
  wire [32:0] r__47;
  wire [31:0] concat_8447;
  wire [32:0] r__45;
  wire [31:0] concat_8369;
  wire [32:0] r__43;
  wire [31:0] concat_8291;
  wire [32:0] r__41;
  wire [31:0] concat_8213;
  wire [32:0] r__39;
  wire [31:0] concat_8135;
  wire [32:0] r__37;
  wire [31:0] concat_8057;
  wire [32:0] r__35;
  wire [31:0] concat_7979;
  wire [32:0] r__33;
  wire [31:0] concat_7901;
  wire [32:0] r__31;
  wire [31:0] concat_7823;
  wire [32:0] r__29;
  wire [31:0] concat_7745;
  wire [32:0] r__27;
  wire [31:0] concat_7667;
  wire [32:0] r__25;
  wire [31:0] concat_7589;
  wire [32:0] r__23;
  wire [31:0] concat_7511;
  wire [32:0] r__21;
  wire [31:0] concat_7433;
  wire [32:0] r__19;
  wire [31:0] concat_7355;
  wire [32:0] r__17;
  wire [31:0] concat_7277;
  wire [32:0] r__15;
  wire [31:0] concat_7199;
  wire [32:0] r__13;
  wire [31:0] concat_7121;
  wire [32:0] r__11;
  wire [31:0] concat_7043;
  wire [32:0] r__9;
  wire [31:0] concat_6965;
  wire [32:0] r__7;
  wire [31:0] concat_6887;
  wire [32:0] r__5;
  wire [31:0] concat_6809;
  wire [32:0] r__3;
  wire [32:0] bivisor__1;
  wire [31:0] concat_6731;
  wire [31:0] concat_6650;
  wire p1_data_enable;
  wire p1_not_valid;
  wire [32:0] r__63;
  wire uge_8994;
  wire [31:0] sub_8995;
  wire uge_8916;
  wire [31:0] sub_8917;
  wire uge_8838;
  wire [31:0] sub_8839;
  wire uge_8760;
  wire [31:0] sub_8761;
  wire uge_8682;
  wire [31:0] sub_8683;
  wire uge_8604;
  wire [31:0] sub_8605;
  wire uge_8526;
  wire [31:0] sub_8527;
  wire uge_8448;
  wire [31:0] sub_8449;
  wire uge_8370;
  wire [31:0] sub_8371;
  wire uge_8292;
  wire [31:0] sub_8293;
  wire uge_8214;
  wire [31:0] sub_8215;
  wire uge_8136;
  wire [31:0] sub_8137;
  wire uge_8058;
  wire [31:0] sub_8059;
  wire uge_7980;
  wire [31:0] sub_7981;
  wire uge_7902;
  wire [31:0] sub_7903;
  wire uge_7824;
  wire [31:0] sub_7825;
  wire uge_7746;
  wire [31:0] sub_7747;
  wire uge_7668;
  wire [31:0] sub_7669;
  wire uge_7590;
  wire [31:0] sub_7591;
  wire uge_7512;
  wire [31:0] sub_7513;
  wire uge_7434;
  wire [31:0] sub_7435;
  wire uge_7356;
  wire [31:0] sub_7357;
  wire uge_7278;
  wire [31:0] sub_7279;
  wire uge_7200;
  wire [31:0] sub_7201;
  wire uge_7122;
  wire [31:0] sub_7123;
  wire uge_7044;
  wire [31:0] sub_7045;
  wire uge_6966;
  wire [31:0] sub_6967;
  wire uge_6888;
  wire [31:0] sub_6889;
  wire uge_6810;
  wire [31:0] sub_6811;
  wire uge_6732;
  wire [31:0] sub_6733;
  wire uge_6652;
  wire [31:0] sub_6653;
  wire p0_enable;
  wire q__32_squeezed_portion_0_width_1;
  wire p34_enable;
  wire p33_enable;
  wire p32_enable;
  wire [31:0] r__62;
  wire [31:0] r__60;
  wire [31:0] r__58;
  wire [31:0] r__56;
  wire [31:0] r__54;
  wire [31:0] r__52;
  wire [31:0] r__50;
  wire [31:0] r__48;
  wire [31:0] r__46;
  wire [31:0] r__44;
  wire [31:0] r__42;
  wire [31:0] r__40;
  wire [31:0] r__38;
  wire [31:0] r__36;
  wire [31:0] r__34;
  wire [31:0] r__32;
  wire [31:0] r__30;
  wire [31:0] r__28;
  wire [31:0] r__26;
  wire [31:0] r__24;
  wire [31:0] r__22;
  wire [31:0] r__20;
  wire [31:0] r__18;
  wire [31:0] r__16;
  wire [31:0] r__14;
  wire [31:0] r__12;
  wire [31:0] r__10;
  wire [31:0] r__8;
  wire [31:0] r__6;
  wire [31:0] r__4;
  wire [31:0] r__2;
  wire bit_slice_6544;
  wire p0_data_enable;
  wire bit_slice_6545;
  wire bit_slice_6546;
  wire bit_slice_6547;
  wire bit_slice_6548;
  wire bit_slice_6549;
  wire bit_slice_6550;
  wire bit_slice_6551;
  wire bit_slice_6552;
  wire bit_slice_6553;
  wire bit_slice_6554;
  wire bit_slice_6555;
  wire bit_slice_6556;
  wire bit_slice_6557;
  wire bit_slice_6558;
  wire bit_slice_6559;
  wire bit_slice_6560;
  wire bit_slice_6561;
  wire bit_slice_6562;
  wire bit_slice_6563;
  wire bit_slice_6564;
  wire bit_slice_6565;
  wire bit_slice_6566;
  wire bit_slice_6567;
  wire bit_slice_6568;
  wire bit_slice_6569;
  wire bit_slice_6570;
  wire bit_slice_6571;
  wire bit_slice_6572;
  wire bit_slice_6573;
  wire bit_slice_6574;
  wire bit_slice_6575;
  wire [31:0] q__32;
  assign xls_float_ips__result_valid_inv = ~__xls_float_ips__result_valid_reg;
  assign xls_float_ips__result_valid_load_en = xls_float_ips__result_rdy | xls_float_ips__result_valid_inv;
  assign xls_float_ips__result_load_en = p31_valid & xls_float_ips__result_valid_load_en;
  assign p32_stage_done = p31_valid & xls_float_ips__result_load_en;
  assign p32_not_valid = ~p31_valid;
  assign p31_enable = p32_stage_done | p32_not_valid;
  assign p31_data_enable = p31_enable & p30_valid;
  assign p31_not_valid = ~p30_valid;
  assign p30_enable = p31_data_enable | p31_not_valid;
  assign p30_data_enable = p30_enable & p29_valid;
  assign p30_not_valid = ~p29_valid;
  assign p29_enable = p30_data_enable | p30_not_valid;
  assign p29_data_enable = p29_enable & p28_valid;
  assign p29_not_valid = ~p28_valid;
  assign p28_enable = p29_data_enable | p29_not_valid;
  assign p28_data_enable = p28_enable & p27_valid;
  assign p28_not_valid = ~p27_valid;
  assign p27_enable = p28_data_enable | p28_not_valid;
  assign p27_data_enable = p27_enable & p26_valid;
  assign p27_not_valid = ~p26_valid;
  assign p26_enable = p27_data_enable | p27_not_valid;
  assign p26_data_enable = p26_enable & p25_valid;
  assign p26_not_valid = ~p25_valid;
  assign p25_enable = p26_data_enable | p26_not_valid;
  assign p25_data_enable = p25_enable & p24_valid;
  assign p25_not_valid = ~p24_valid;
  assign p24_enable = p25_data_enable | p25_not_valid;
  assign p24_data_enable = p24_enable & p23_valid;
  assign p24_not_valid = ~p23_valid;
  assign p23_enable = p24_data_enable | p24_not_valid;
  assign p23_data_enable = p23_enable & p22_valid;
  assign p23_not_valid = ~p22_valid;
  assign p22_enable = p23_data_enable | p23_not_valid;
  assign p22_data_enable = p22_enable & p21_valid;
  assign p22_not_valid = ~p21_valid;
  assign p21_enable = p22_data_enable | p22_not_valid;
  assign p21_data_enable = p21_enable & p20_valid;
  assign p21_not_valid = ~p20_valid;
  assign p20_enable = p21_data_enable | p21_not_valid;
  assign p20_data_enable = p20_enable & p19_valid;
  assign p20_not_valid = ~p19_valid;
  assign p19_enable = p20_data_enable | p20_not_valid;
  assign p19_data_enable = p19_enable & p18_valid;
  assign p19_not_valid = ~p18_valid;
  assign p18_enable = p19_data_enable | p19_not_valid;
  assign p18_data_enable = p18_enable & p17_valid;
  assign p18_not_valid = ~p17_valid;
  assign p17_enable = p18_data_enable | p18_not_valid;
  assign p17_data_enable = p17_enable & p16_valid;
  assign p17_not_valid = ~p16_valid;
  assign p16_enable = p17_data_enable | p17_not_valid;
  assign p16_data_enable = p16_enable & p15_valid;
  assign p16_not_valid = ~p15_valid;
  assign p15_enable = p16_data_enable | p16_not_valid;
  assign p15_data_enable = p15_enable & p14_valid;
  assign p15_not_valid = ~p14_valid;
  assign p14_enable = p15_data_enable | p15_not_valid;
  assign p14_data_enable = p14_enable & p13_valid;
  assign p14_not_valid = ~p13_valid;
  assign p13_enable = p14_data_enable | p14_not_valid;
  assign p13_data_enable = p13_enable & p12_valid;
  assign p13_not_valid = ~p12_valid;
  assign p12_enable = p13_data_enable | p13_not_valid;
  assign p12_data_enable = p12_enable & p11_valid;
  assign p12_not_valid = ~p11_valid;
  assign p11_enable = p12_data_enable | p12_not_valid;
  assign p11_data_enable = p11_enable & p10_valid;
  assign p11_not_valid = ~p10_valid;
  assign p10_enable = p11_data_enable | p11_not_valid;
  assign p10_data_enable = p10_enable & p9_valid;
  assign p10_not_valid = ~p9_valid;
  assign p9_enable = p10_data_enable | p10_not_valid;
  assign p9_data_enable = p9_enable & p8_valid;
  assign p9_not_valid = ~p8_valid;
  assign p8_enable = p9_data_enable | p9_not_valid;
  assign p8_data_enable = p8_enable & p7_valid;
  assign p8_not_valid = ~p7_valid;
  assign p7_enable = p8_data_enable | p8_not_valid;
  assign p7_data_enable = p7_enable & p6_valid;
  assign p7_not_valid = ~p6_valid;
  assign p6_enable = p7_data_enable | p7_not_valid;
  assign p6_data_enable = p6_enable & p5_valid;
  assign p6_not_valid = ~p5_valid;
  assign p5_enable = p6_data_enable | p6_not_valid;
  assign p5_data_enable = p5_enable & p4_valid;
  assign p5_not_valid = ~p4_valid;
  assign p4_enable = p5_data_enable | p5_not_valid;
  assign p4_data_enable = p4_enable & p3_valid;
  assign p4_not_valid = ~p3_valid;
  assign p3_enable = p4_data_enable | p4_not_valid;
  assign p3_data_enable = p3_enable & p2_valid;
  assign p3_not_valid = ~p2_valid;
  assign p2_enable = p3_data_enable | p3_not_valid;
  assign p2_data_enable = p2_enable & p1_valid;
  assign p2_not_valid = ~p1_valid;
  assign p1_enable = p2_data_enable | p2_not_valid;
  assign p1_stage_done = p0_valid & xls_float_ips__rhs_vld;
  assign r__61 = {p30_r__60, p30_bit_slice_6574};
  assign concat_8993 = {p30_r__60[30:0], p30_bit_slice_6574};
  assign r__59 = {p29_r__58, p29_bit_slice_6573};
  assign concat_8915 = {p29_r__58[30:0], p29_bit_slice_6573};
  assign r__57 = {p28_r__56, p28_bit_slice_6572};
  assign concat_8837 = {p28_r__56[30:0], p28_bit_slice_6572};
  assign r__55 = {p27_r__54, p27_bit_slice_6571};
  assign concat_8759 = {p27_r__54[30:0], p27_bit_slice_6571};
  assign r__53 = {p26_r__52, p26_bit_slice_6570};
  assign concat_8681 = {p26_r__52[30:0], p26_bit_slice_6570};
  assign r__51 = {p25_r__50, p25_bit_slice_6569};
  assign concat_8603 = {p25_r__50[30:0], p25_bit_slice_6569};
  assign r__49 = {p24_r__48, p24_bit_slice_6568};
  assign concat_8525 = {p24_r__48[30:0], p24_bit_slice_6568};
  assign r__47 = {p23_r__46, p23_bit_slice_6567};
  assign concat_8447 = {p23_r__46[30:0], p23_bit_slice_6567};
  assign r__45 = {p22_r__44, p22_bit_slice_6566};
  assign concat_8369 = {p22_r__44[30:0], p22_bit_slice_6566};
  assign r__43 = {p21_r__42, p21_bit_slice_6565};
  assign concat_8291 = {p21_r__42[30:0], p21_bit_slice_6565};
  assign r__41 = {p20_r__40, p20_bit_slice_6564};
  assign concat_8213 = {p20_r__40[30:0], p20_bit_slice_6564};
  assign r__39 = {p19_r__38, p19_bit_slice_6563};
  assign concat_8135 = {p19_r__38[30:0], p19_bit_slice_6563};
  assign r__37 = {p18_r__36, p18_bit_slice_6562};
  assign concat_8057 = {p18_r__36[30:0], p18_bit_slice_6562};
  assign r__35 = {p17_r__34, p17_bit_slice_6561};
  assign concat_7979 = {p17_r__34[30:0], p17_bit_slice_6561};
  assign r__33 = {p16_r__32, p16_bit_slice_6560};
  assign concat_7901 = {p16_r__32[30:0], p16_bit_slice_6560};
  assign r__31 = {p15_r__30, p15_bit_slice_6559};
  assign concat_7823 = {p15_r__30[30:0], p15_bit_slice_6559};
  assign r__29 = {p14_r__28, p14_bit_slice_6558};
  assign concat_7745 = {p14_r__28[30:0], p14_bit_slice_6558};
  assign r__27 = {p13_r__26, p13_bit_slice_6557};
  assign concat_7667 = {p13_r__26[30:0], p13_bit_slice_6557};
  assign r__25 = {p12_r__24, p12_bit_slice_6556};
  assign concat_7589 = {p12_r__24[30:0], p12_bit_slice_6556};
  assign r__23 = {p11_r__22, p11_bit_slice_6555};
  assign concat_7511 = {p11_r__22[30:0], p11_bit_slice_6555};
  assign r__21 = {p10_r__20, p10_bit_slice_6554};
  assign concat_7433 = {p10_r__20[30:0], p10_bit_slice_6554};
  assign r__19 = {p9_r__18, p9_bit_slice_6553};
  assign concat_7355 = {p9_r__18[30:0], p9_bit_slice_6553};
  assign r__17 = {p8_r__16, p8_bit_slice_6552};
  assign concat_7277 = {p8_r__16[30:0], p8_bit_slice_6552};
  assign r__15 = {p7_r__14, p7_bit_slice_6551};
  assign concat_7199 = {p7_r__14[30:0], p7_bit_slice_6551};
  assign r__13 = {p6_r__12, p6_bit_slice_6550};
  assign concat_7121 = {p6_r__12[30:0], p6_bit_slice_6550};
  assign r__11 = {p5_r__10, p5_bit_slice_6549};
  assign concat_7043 = {p5_r__10[30:0], p5_bit_slice_6549};
  assign r__9 = {p4_r__8, p4_bit_slice_6548};
  assign concat_6965 = {p4_r__8[30:0], p4_bit_slice_6548};
  assign r__7 = {p3_r__6, p3_bit_slice_6547};
  assign concat_6887 = {p3_r__6[30:0], p3_bit_slice_6547};
  assign r__5 = {p2_r__4, p2_bit_slice_6546};
  assign concat_6809 = {p2_r__4[30:0], p2_bit_slice_6546};
  assign r__3 = {p1_r__2, p1_bit_slice_6545};
  assign bivisor__1 = {1'h0, p1_b};
  assign concat_6731 = {p1_r__2[30:0], p1_bit_slice_6545};
  assign concat_6650 = {31'h0000_0000, p0_bit_slice_6544};
  assign p1_data_enable = p1_enable & p1_stage_done;
  assign p1_not_valid = ~p0_valid;
  assign r__63 = {p31_r__62, p31_bit_slice_6575};
  assign uge_8994 = r__61 >= p30_bivisor__1;
  assign sub_8995 = concat_8993 - p30_b;
  assign uge_8916 = r__59 >= p29_bivisor__1;
  assign sub_8917 = concat_8915 - p29_b;
  assign uge_8838 = r__57 >= p28_bivisor__1;
  assign sub_8839 = concat_8837 - p28_b;
  assign uge_8760 = r__55 >= p27_bivisor__1;
  assign sub_8761 = concat_8759 - p27_b;
  assign uge_8682 = r__53 >= p26_bivisor__1;
  assign sub_8683 = concat_8681 - p26_b;
  assign uge_8604 = r__51 >= p25_bivisor__1;
  assign sub_8605 = concat_8603 - p25_b;
  assign uge_8526 = r__49 >= p24_bivisor__1;
  assign sub_8527 = concat_8525 - p24_b;
  assign uge_8448 = r__47 >= p23_bivisor__1;
  assign sub_8449 = concat_8447 - p23_b;
  assign uge_8370 = r__45 >= p22_bivisor__1;
  assign sub_8371 = concat_8369 - p22_b;
  assign uge_8292 = r__43 >= p21_bivisor__1;
  assign sub_8293 = concat_8291 - p21_b;
  assign uge_8214 = r__41 >= p20_bivisor__1;
  assign sub_8215 = concat_8213 - p20_b;
  assign uge_8136 = r__39 >= p19_bivisor__1;
  assign sub_8137 = concat_8135 - p19_b;
  assign uge_8058 = r__37 >= p18_bivisor__1;
  assign sub_8059 = concat_8057 - p18_b;
  assign uge_7980 = r__35 >= p17_bivisor__1;
  assign sub_7981 = concat_7979 - p17_b;
  assign uge_7902 = r__33 >= p16_bivisor__1;
  assign sub_7903 = concat_7901 - p16_b;
  assign uge_7824 = r__31 >= p15_bivisor__1;
  assign sub_7825 = concat_7823 - p15_b;
  assign uge_7746 = r__29 >= p14_bivisor__1;
  assign sub_7747 = concat_7745 - p14_b;
  assign uge_7668 = r__27 >= p13_bivisor__1;
  assign sub_7669 = concat_7667 - p13_b;
  assign uge_7590 = r__25 >= p12_bivisor__1;
  assign sub_7591 = concat_7589 - p12_b;
  assign uge_7512 = r__23 >= p11_bivisor__1;
  assign sub_7513 = concat_7511 - p11_b;
  assign uge_7434 = r__21 >= p10_bivisor__1;
  assign sub_7435 = concat_7433 - p10_b;
  assign uge_7356 = r__19 >= p9_bivisor__1;
  assign sub_7357 = concat_7355 - p9_b;
  assign uge_7278 = r__17 >= p8_bivisor__1;
  assign sub_7279 = concat_7277 - p8_b;
  assign uge_7200 = r__15 >= p7_bivisor__1;
  assign sub_7201 = concat_7199 - p7_b;
  assign uge_7122 = r__13 >= p6_bivisor__1;
  assign sub_7123 = concat_7121 - p6_b;
  assign uge_7044 = r__11 >= p5_bivisor__1;
  assign sub_7045 = concat_7043 - p5_b;
  assign uge_6966 = r__9 >= p4_bivisor__1;
  assign sub_6967 = concat_6965 - p4_b;
  assign uge_6888 = r__7 >= p3_bivisor__1;
  assign sub_6889 = concat_6887 - p3_b;
  assign uge_6810 = r__5 >= p2_bivisor__1;
  assign sub_6811 = concat_6809 - p2_b;
  assign uge_6732 = r__3 >= bivisor__1;
  assign sub_6733 = concat_6731 - p1_b;
  assign uge_6652 = concat_6650 >= xls_float_ips__rhs;
  assign sub_6653 = concat_6650 - xls_float_ips__rhs;
  assign p0_enable = p1_data_enable | p1_not_valid;
  assign q__32_squeezed_portion_0_width_1 = r__63 >= p31_bivisor__1;
  assign p34_enable = 1'h1;
  assign p33_enable = 1'h1;
  assign p32_enable = 1'h1;
  assign r__62 = uge_8994 ? sub_8995 : concat_8993;
  assign r__60 = uge_8916 ? sub_8917 : concat_8915;
  assign r__58 = uge_8838 ? sub_8839 : concat_8837;
  assign r__56 = uge_8760 ? sub_8761 : concat_8759;
  assign r__54 = uge_8682 ? sub_8683 : concat_8681;
  assign r__52 = uge_8604 ? sub_8605 : concat_8603;
  assign r__50 = uge_8526 ? sub_8527 : concat_8525;
  assign r__48 = uge_8448 ? sub_8449 : concat_8447;
  assign r__46 = uge_8370 ? sub_8371 : concat_8369;
  assign r__44 = uge_8292 ? sub_8293 : concat_8291;
  assign r__42 = uge_8214 ? sub_8215 : concat_8213;
  assign r__40 = uge_8136 ? sub_8137 : concat_8135;
  assign r__38 = uge_8058 ? sub_8059 : concat_8057;
  assign r__36 = uge_7980 ? sub_7981 : concat_7979;
  assign r__34 = uge_7902 ? sub_7903 : concat_7901;
  assign r__32 = uge_7824 ? sub_7825 : concat_7823;
  assign r__30 = uge_7746 ? sub_7747 : concat_7745;
  assign r__28 = uge_7668 ? sub_7669 : concat_7667;
  assign r__26 = uge_7590 ? sub_7591 : concat_7589;
  assign r__24 = uge_7512 ? sub_7513 : concat_7511;
  assign r__22 = uge_7434 ? sub_7435 : concat_7433;
  assign r__20 = uge_7356 ? sub_7357 : concat_7355;
  assign r__18 = uge_7278 ? sub_7279 : concat_7277;
  assign r__16 = uge_7200 ? sub_7201 : concat_7199;
  assign r__14 = uge_7122 ? sub_7123 : concat_7121;
  assign r__12 = uge_7044 ? sub_7045 : concat_7043;
  assign r__10 = uge_6966 ? sub_6967 : concat_6965;
  assign r__8 = uge_6888 ? sub_6889 : concat_6887;
  assign r__6 = uge_6810 ? sub_6811 : concat_6809;
  assign r__4 = uge_6732 ? sub_6733 : concat_6731;
  assign r__2 = uge_6652 ? sub_6653 : concat_6650;
  assign bit_slice_6544 = xls_float_ips__lhs[31];
  assign p0_data_enable = p0_enable & xls_float_ips__lhs_vld;
  assign bit_slice_6545 = xls_float_ips__lhs[30];
  assign bit_slice_6546 = xls_float_ips__lhs[29];
  assign bit_slice_6547 = xls_float_ips__lhs[28];
  assign bit_slice_6548 = xls_float_ips__lhs[27];
  assign bit_slice_6549 = xls_float_ips__lhs[26];
  assign bit_slice_6550 = xls_float_ips__lhs[25];
  assign bit_slice_6551 = xls_float_ips__lhs[24];
  assign bit_slice_6552 = xls_float_ips__lhs[23];
  assign bit_slice_6553 = xls_float_ips__lhs[22];
  assign bit_slice_6554 = xls_float_ips__lhs[21];
  assign bit_slice_6555 = xls_float_ips__lhs[20];
  assign bit_slice_6556 = xls_float_ips__lhs[19];
  assign bit_slice_6557 = xls_float_ips__lhs[18];
  assign bit_slice_6558 = xls_float_ips__lhs[17];
  assign bit_slice_6559 = xls_float_ips__lhs[16];
  assign bit_slice_6560 = xls_float_ips__lhs[15];
  assign bit_slice_6561 = xls_float_ips__lhs[14];
  assign bit_slice_6562 = xls_float_ips__lhs[13];
  assign bit_slice_6563 = xls_float_ips__lhs[12];
  assign bit_slice_6564 = xls_float_ips__lhs[11];
  assign bit_slice_6565 = xls_float_ips__lhs[10];
  assign bit_slice_6566 = xls_float_ips__lhs[9];
  assign bit_slice_6567 = xls_float_ips__lhs[8];
  assign bit_slice_6568 = xls_float_ips__lhs[7];
  assign bit_slice_6569 = xls_float_ips__lhs[6];
  assign bit_slice_6570 = xls_float_ips__lhs[5];
  assign bit_slice_6571 = xls_float_ips__lhs[4];
  assign bit_slice_6572 = xls_float_ips__lhs[3];
  assign bit_slice_6573 = xls_float_ips__lhs[2];
  assign bit_slice_6574 = xls_float_ips__lhs[1];
  assign bit_slice_6575 = xls_float_ips__lhs[0];
  assign q__32 = {p31_uge_6652, p31_uge_6732, p31_uge_6810, p31_uge_6888, p31_uge_6966, p31_uge_7044, p31_uge_7122, p31_uge_7200, p31_uge_7278, p31_uge_7356, p31_uge_7434, p31_uge_7512, p31_uge_7590, p31_uge_7668, p31_uge_7746, p31_uge_7824, p31_uge_7902, p31_uge_7980, p31_uge_8058, p31_uge_8136, p31_uge_8214, p31_uge_8292, p31_uge_8370, p31_uge_8448, p31_uge_8526, p31_uge_8604, p31_uge_8682, p31_uge_8760, p31_uge_8838, p31_uge_8916, p31_uge_8994, q__32_squeezed_portion_0_width_1};
  always @ (posedge clk) begin
    if (rst) begin
      p0_bit_slice_6544 <= 1'h0;
      p0_bit_slice_6545 <= 1'h0;
      p0_bit_slice_6546 <= 1'h0;
      p0_bit_slice_6547 <= 1'h0;
      p0_bit_slice_6548 <= 1'h0;
      p0_bit_slice_6549 <= 1'h0;
      p0_bit_slice_6550 <= 1'h0;
      p0_bit_slice_6551 <= 1'h0;
      p0_bit_slice_6552 <= 1'h0;
      p0_bit_slice_6553 <= 1'h0;
      p0_bit_slice_6554 <= 1'h0;
      p0_bit_slice_6555 <= 1'h0;
      p0_bit_slice_6556 <= 1'h0;
      p0_bit_slice_6557 <= 1'h0;
      p0_bit_slice_6558 <= 1'h0;
      p0_bit_slice_6559 <= 1'h0;
      p0_bit_slice_6560 <= 1'h0;
      p0_bit_slice_6561 <= 1'h0;
      p0_bit_slice_6562 <= 1'h0;
      p0_bit_slice_6563 <= 1'h0;
      p0_bit_slice_6564 <= 1'h0;
      p0_bit_slice_6565 <= 1'h0;
      p0_bit_slice_6566 <= 1'h0;
      p0_bit_slice_6567 <= 1'h0;
      p0_bit_slice_6568 <= 1'h0;
      p0_bit_slice_6569 <= 1'h0;
      p0_bit_slice_6570 <= 1'h0;
      p0_bit_slice_6571 <= 1'h0;
      p0_bit_slice_6572 <= 1'h0;
      p0_bit_slice_6573 <= 1'h0;
      p0_bit_slice_6574 <= 1'h0;
      p0_bit_slice_6575 <= 1'h0;
      p1_b <= 32'h0000_0000;
      p1_uge_6652 <= 1'h0;
      p1_r__2 <= 32'h0000_0000;
      p1_bit_slice_6545 <= 1'h0;
      p1_bit_slice_6546 <= 1'h0;
      p1_bit_slice_6547 <= 1'h0;
      p1_bit_slice_6548 <= 1'h0;
      p1_bit_slice_6549 <= 1'h0;
      p1_bit_slice_6550 <= 1'h0;
      p1_bit_slice_6551 <= 1'h0;
      p1_bit_slice_6552 <= 1'h0;
      p1_bit_slice_6553 <= 1'h0;
      p1_bit_slice_6554 <= 1'h0;
      p1_bit_slice_6555 <= 1'h0;
      p1_bit_slice_6556 <= 1'h0;
      p1_bit_slice_6557 <= 1'h0;
      p1_bit_slice_6558 <= 1'h0;
      p1_bit_slice_6559 <= 1'h0;
      p1_bit_slice_6560 <= 1'h0;
      p1_bit_slice_6561 <= 1'h0;
      p1_bit_slice_6562 <= 1'h0;
      p1_bit_slice_6563 <= 1'h0;
      p1_bit_slice_6564 <= 1'h0;
      p1_bit_slice_6565 <= 1'h0;
      p1_bit_slice_6566 <= 1'h0;
      p1_bit_slice_6567 <= 1'h0;
      p1_bit_slice_6568 <= 1'h0;
      p1_bit_slice_6569 <= 1'h0;
      p1_bit_slice_6570 <= 1'h0;
      p1_bit_slice_6571 <= 1'h0;
      p1_bit_slice_6572 <= 1'h0;
      p1_bit_slice_6573 <= 1'h0;
      p1_bit_slice_6574 <= 1'h0;
      p1_bit_slice_6575 <= 1'h0;
      p2_b <= 32'h0000_0000;
      p2_uge_6652 <= 1'h0;
      p2_bivisor__1 <= 33'h0_0000_0000;
      p2_uge_6732 <= 1'h0;
      p2_r__4 <= 32'h0000_0000;
      p2_bit_slice_6546 <= 1'h0;
      p2_bit_slice_6547 <= 1'h0;
      p2_bit_slice_6548 <= 1'h0;
      p2_bit_slice_6549 <= 1'h0;
      p2_bit_slice_6550 <= 1'h0;
      p2_bit_slice_6551 <= 1'h0;
      p2_bit_slice_6552 <= 1'h0;
      p2_bit_slice_6553 <= 1'h0;
      p2_bit_slice_6554 <= 1'h0;
      p2_bit_slice_6555 <= 1'h0;
      p2_bit_slice_6556 <= 1'h0;
      p2_bit_slice_6557 <= 1'h0;
      p2_bit_slice_6558 <= 1'h0;
      p2_bit_slice_6559 <= 1'h0;
      p2_bit_slice_6560 <= 1'h0;
      p2_bit_slice_6561 <= 1'h0;
      p2_bit_slice_6562 <= 1'h0;
      p2_bit_slice_6563 <= 1'h0;
      p2_bit_slice_6564 <= 1'h0;
      p2_bit_slice_6565 <= 1'h0;
      p2_bit_slice_6566 <= 1'h0;
      p2_bit_slice_6567 <= 1'h0;
      p2_bit_slice_6568 <= 1'h0;
      p2_bit_slice_6569 <= 1'h0;
      p2_bit_slice_6570 <= 1'h0;
      p2_bit_slice_6571 <= 1'h0;
      p2_bit_slice_6572 <= 1'h0;
      p2_bit_slice_6573 <= 1'h0;
      p2_bit_slice_6574 <= 1'h0;
      p2_bit_slice_6575 <= 1'h0;
      p3_b <= 32'h0000_0000;
      p3_uge_6652 <= 1'h0;
      p3_bivisor__1 <= 33'h0_0000_0000;
      p3_uge_6732 <= 1'h0;
      p3_uge_6810 <= 1'h0;
      p3_r__6 <= 32'h0000_0000;
      p3_bit_slice_6547 <= 1'h0;
      p3_bit_slice_6548 <= 1'h0;
      p3_bit_slice_6549 <= 1'h0;
      p3_bit_slice_6550 <= 1'h0;
      p3_bit_slice_6551 <= 1'h0;
      p3_bit_slice_6552 <= 1'h0;
      p3_bit_slice_6553 <= 1'h0;
      p3_bit_slice_6554 <= 1'h0;
      p3_bit_slice_6555 <= 1'h0;
      p3_bit_slice_6556 <= 1'h0;
      p3_bit_slice_6557 <= 1'h0;
      p3_bit_slice_6558 <= 1'h0;
      p3_bit_slice_6559 <= 1'h0;
      p3_bit_slice_6560 <= 1'h0;
      p3_bit_slice_6561 <= 1'h0;
      p3_bit_slice_6562 <= 1'h0;
      p3_bit_slice_6563 <= 1'h0;
      p3_bit_slice_6564 <= 1'h0;
      p3_bit_slice_6565 <= 1'h0;
      p3_bit_slice_6566 <= 1'h0;
      p3_bit_slice_6567 <= 1'h0;
      p3_bit_slice_6568 <= 1'h0;
      p3_bit_slice_6569 <= 1'h0;
      p3_bit_slice_6570 <= 1'h0;
      p3_bit_slice_6571 <= 1'h0;
      p3_bit_slice_6572 <= 1'h0;
      p3_bit_slice_6573 <= 1'h0;
      p3_bit_slice_6574 <= 1'h0;
      p3_bit_slice_6575 <= 1'h0;
      p4_b <= 32'h0000_0000;
      p4_uge_6652 <= 1'h0;
      p4_bivisor__1 <= 33'h0_0000_0000;
      p4_uge_6732 <= 1'h0;
      p4_uge_6810 <= 1'h0;
      p4_uge_6888 <= 1'h0;
      p4_r__8 <= 32'h0000_0000;
      p4_bit_slice_6548 <= 1'h0;
      p4_bit_slice_6549 <= 1'h0;
      p4_bit_slice_6550 <= 1'h0;
      p4_bit_slice_6551 <= 1'h0;
      p4_bit_slice_6552 <= 1'h0;
      p4_bit_slice_6553 <= 1'h0;
      p4_bit_slice_6554 <= 1'h0;
      p4_bit_slice_6555 <= 1'h0;
      p4_bit_slice_6556 <= 1'h0;
      p4_bit_slice_6557 <= 1'h0;
      p4_bit_slice_6558 <= 1'h0;
      p4_bit_slice_6559 <= 1'h0;
      p4_bit_slice_6560 <= 1'h0;
      p4_bit_slice_6561 <= 1'h0;
      p4_bit_slice_6562 <= 1'h0;
      p4_bit_slice_6563 <= 1'h0;
      p4_bit_slice_6564 <= 1'h0;
      p4_bit_slice_6565 <= 1'h0;
      p4_bit_slice_6566 <= 1'h0;
      p4_bit_slice_6567 <= 1'h0;
      p4_bit_slice_6568 <= 1'h0;
      p4_bit_slice_6569 <= 1'h0;
      p4_bit_slice_6570 <= 1'h0;
      p4_bit_slice_6571 <= 1'h0;
      p4_bit_slice_6572 <= 1'h0;
      p4_bit_slice_6573 <= 1'h0;
      p4_bit_slice_6574 <= 1'h0;
      p4_bit_slice_6575 <= 1'h0;
      p5_b <= 32'h0000_0000;
      p5_uge_6652 <= 1'h0;
      p5_bivisor__1 <= 33'h0_0000_0000;
      p5_uge_6732 <= 1'h0;
      p5_uge_6810 <= 1'h0;
      p5_uge_6888 <= 1'h0;
      p5_uge_6966 <= 1'h0;
      p5_r__10 <= 32'h0000_0000;
      p5_bit_slice_6549 <= 1'h0;
      p5_bit_slice_6550 <= 1'h0;
      p5_bit_slice_6551 <= 1'h0;
      p5_bit_slice_6552 <= 1'h0;
      p5_bit_slice_6553 <= 1'h0;
      p5_bit_slice_6554 <= 1'h0;
      p5_bit_slice_6555 <= 1'h0;
      p5_bit_slice_6556 <= 1'h0;
      p5_bit_slice_6557 <= 1'h0;
      p5_bit_slice_6558 <= 1'h0;
      p5_bit_slice_6559 <= 1'h0;
      p5_bit_slice_6560 <= 1'h0;
      p5_bit_slice_6561 <= 1'h0;
      p5_bit_slice_6562 <= 1'h0;
      p5_bit_slice_6563 <= 1'h0;
      p5_bit_slice_6564 <= 1'h0;
      p5_bit_slice_6565 <= 1'h0;
      p5_bit_slice_6566 <= 1'h0;
      p5_bit_slice_6567 <= 1'h0;
      p5_bit_slice_6568 <= 1'h0;
      p5_bit_slice_6569 <= 1'h0;
      p5_bit_slice_6570 <= 1'h0;
      p5_bit_slice_6571 <= 1'h0;
      p5_bit_slice_6572 <= 1'h0;
      p5_bit_slice_6573 <= 1'h0;
      p5_bit_slice_6574 <= 1'h0;
      p5_bit_slice_6575 <= 1'h0;
      p6_b <= 32'h0000_0000;
      p6_uge_6652 <= 1'h0;
      p6_bivisor__1 <= 33'h0_0000_0000;
      p6_uge_6732 <= 1'h0;
      p6_uge_6810 <= 1'h0;
      p6_uge_6888 <= 1'h0;
      p6_uge_6966 <= 1'h0;
      p6_uge_7044 <= 1'h0;
      p6_r__12 <= 32'h0000_0000;
      p6_bit_slice_6550 <= 1'h0;
      p6_bit_slice_6551 <= 1'h0;
      p6_bit_slice_6552 <= 1'h0;
      p6_bit_slice_6553 <= 1'h0;
      p6_bit_slice_6554 <= 1'h0;
      p6_bit_slice_6555 <= 1'h0;
      p6_bit_slice_6556 <= 1'h0;
      p6_bit_slice_6557 <= 1'h0;
      p6_bit_slice_6558 <= 1'h0;
      p6_bit_slice_6559 <= 1'h0;
      p6_bit_slice_6560 <= 1'h0;
      p6_bit_slice_6561 <= 1'h0;
      p6_bit_slice_6562 <= 1'h0;
      p6_bit_slice_6563 <= 1'h0;
      p6_bit_slice_6564 <= 1'h0;
      p6_bit_slice_6565 <= 1'h0;
      p6_bit_slice_6566 <= 1'h0;
      p6_bit_slice_6567 <= 1'h0;
      p6_bit_slice_6568 <= 1'h0;
      p6_bit_slice_6569 <= 1'h0;
      p6_bit_slice_6570 <= 1'h0;
      p6_bit_slice_6571 <= 1'h0;
      p6_bit_slice_6572 <= 1'h0;
      p6_bit_slice_6573 <= 1'h0;
      p6_bit_slice_6574 <= 1'h0;
      p6_bit_slice_6575 <= 1'h0;
      p7_b <= 32'h0000_0000;
      p7_uge_6652 <= 1'h0;
      p7_bivisor__1 <= 33'h0_0000_0000;
      p7_uge_6732 <= 1'h0;
      p7_uge_6810 <= 1'h0;
      p7_uge_6888 <= 1'h0;
      p7_uge_6966 <= 1'h0;
      p7_uge_7044 <= 1'h0;
      p7_uge_7122 <= 1'h0;
      p7_r__14 <= 32'h0000_0000;
      p7_bit_slice_6551 <= 1'h0;
      p7_bit_slice_6552 <= 1'h0;
      p7_bit_slice_6553 <= 1'h0;
      p7_bit_slice_6554 <= 1'h0;
      p7_bit_slice_6555 <= 1'h0;
      p7_bit_slice_6556 <= 1'h0;
      p7_bit_slice_6557 <= 1'h0;
      p7_bit_slice_6558 <= 1'h0;
      p7_bit_slice_6559 <= 1'h0;
      p7_bit_slice_6560 <= 1'h0;
      p7_bit_slice_6561 <= 1'h0;
      p7_bit_slice_6562 <= 1'h0;
      p7_bit_slice_6563 <= 1'h0;
      p7_bit_slice_6564 <= 1'h0;
      p7_bit_slice_6565 <= 1'h0;
      p7_bit_slice_6566 <= 1'h0;
      p7_bit_slice_6567 <= 1'h0;
      p7_bit_slice_6568 <= 1'h0;
      p7_bit_slice_6569 <= 1'h0;
      p7_bit_slice_6570 <= 1'h0;
      p7_bit_slice_6571 <= 1'h0;
      p7_bit_slice_6572 <= 1'h0;
      p7_bit_slice_6573 <= 1'h0;
      p7_bit_slice_6574 <= 1'h0;
      p7_bit_slice_6575 <= 1'h0;
      p8_b <= 32'h0000_0000;
      p8_uge_6652 <= 1'h0;
      p8_bivisor__1 <= 33'h0_0000_0000;
      p8_uge_6732 <= 1'h0;
      p8_uge_6810 <= 1'h0;
      p8_uge_6888 <= 1'h0;
      p8_uge_6966 <= 1'h0;
      p8_uge_7044 <= 1'h0;
      p8_uge_7122 <= 1'h0;
      p8_uge_7200 <= 1'h0;
      p8_r__16 <= 32'h0000_0000;
      p8_bit_slice_6552 <= 1'h0;
      p8_bit_slice_6553 <= 1'h0;
      p8_bit_slice_6554 <= 1'h0;
      p8_bit_slice_6555 <= 1'h0;
      p8_bit_slice_6556 <= 1'h0;
      p8_bit_slice_6557 <= 1'h0;
      p8_bit_slice_6558 <= 1'h0;
      p8_bit_slice_6559 <= 1'h0;
      p8_bit_slice_6560 <= 1'h0;
      p8_bit_slice_6561 <= 1'h0;
      p8_bit_slice_6562 <= 1'h0;
      p8_bit_slice_6563 <= 1'h0;
      p8_bit_slice_6564 <= 1'h0;
      p8_bit_slice_6565 <= 1'h0;
      p8_bit_slice_6566 <= 1'h0;
      p8_bit_slice_6567 <= 1'h0;
      p8_bit_slice_6568 <= 1'h0;
      p8_bit_slice_6569 <= 1'h0;
      p8_bit_slice_6570 <= 1'h0;
      p8_bit_slice_6571 <= 1'h0;
      p8_bit_slice_6572 <= 1'h0;
      p8_bit_slice_6573 <= 1'h0;
      p8_bit_slice_6574 <= 1'h0;
      p8_bit_slice_6575 <= 1'h0;
      p9_b <= 32'h0000_0000;
      p9_uge_6652 <= 1'h0;
      p9_bivisor__1 <= 33'h0_0000_0000;
      p9_uge_6732 <= 1'h0;
      p9_uge_6810 <= 1'h0;
      p9_uge_6888 <= 1'h0;
      p9_uge_6966 <= 1'h0;
      p9_uge_7044 <= 1'h0;
      p9_uge_7122 <= 1'h0;
      p9_uge_7200 <= 1'h0;
      p9_uge_7278 <= 1'h0;
      p9_r__18 <= 32'h0000_0000;
      p9_bit_slice_6553 <= 1'h0;
      p9_bit_slice_6554 <= 1'h0;
      p9_bit_slice_6555 <= 1'h0;
      p9_bit_slice_6556 <= 1'h0;
      p9_bit_slice_6557 <= 1'h0;
      p9_bit_slice_6558 <= 1'h0;
      p9_bit_slice_6559 <= 1'h0;
      p9_bit_slice_6560 <= 1'h0;
      p9_bit_slice_6561 <= 1'h0;
      p9_bit_slice_6562 <= 1'h0;
      p9_bit_slice_6563 <= 1'h0;
      p9_bit_slice_6564 <= 1'h0;
      p9_bit_slice_6565 <= 1'h0;
      p9_bit_slice_6566 <= 1'h0;
      p9_bit_slice_6567 <= 1'h0;
      p9_bit_slice_6568 <= 1'h0;
      p9_bit_slice_6569 <= 1'h0;
      p9_bit_slice_6570 <= 1'h0;
      p9_bit_slice_6571 <= 1'h0;
      p9_bit_slice_6572 <= 1'h0;
      p9_bit_slice_6573 <= 1'h0;
      p9_bit_slice_6574 <= 1'h0;
      p9_bit_slice_6575 <= 1'h0;
      p10_b <= 32'h0000_0000;
      p10_uge_6652 <= 1'h0;
      p10_bivisor__1 <= 33'h0_0000_0000;
      p10_uge_6732 <= 1'h0;
      p10_uge_6810 <= 1'h0;
      p10_uge_6888 <= 1'h0;
      p10_uge_6966 <= 1'h0;
      p10_uge_7044 <= 1'h0;
      p10_uge_7122 <= 1'h0;
      p10_uge_7200 <= 1'h0;
      p10_uge_7278 <= 1'h0;
      p10_uge_7356 <= 1'h0;
      p10_r__20 <= 32'h0000_0000;
      p10_bit_slice_6554 <= 1'h0;
      p10_bit_slice_6555 <= 1'h0;
      p10_bit_slice_6556 <= 1'h0;
      p10_bit_slice_6557 <= 1'h0;
      p10_bit_slice_6558 <= 1'h0;
      p10_bit_slice_6559 <= 1'h0;
      p10_bit_slice_6560 <= 1'h0;
      p10_bit_slice_6561 <= 1'h0;
      p10_bit_slice_6562 <= 1'h0;
      p10_bit_slice_6563 <= 1'h0;
      p10_bit_slice_6564 <= 1'h0;
      p10_bit_slice_6565 <= 1'h0;
      p10_bit_slice_6566 <= 1'h0;
      p10_bit_slice_6567 <= 1'h0;
      p10_bit_slice_6568 <= 1'h0;
      p10_bit_slice_6569 <= 1'h0;
      p10_bit_slice_6570 <= 1'h0;
      p10_bit_slice_6571 <= 1'h0;
      p10_bit_slice_6572 <= 1'h0;
      p10_bit_slice_6573 <= 1'h0;
      p10_bit_slice_6574 <= 1'h0;
      p10_bit_slice_6575 <= 1'h0;
      p11_b <= 32'h0000_0000;
      p11_uge_6652 <= 1'h0;
      p11_bivisor__1 <= 33'h0_0000_0000;
      p11_uge_6732 <= 1'h0;
      p11_uge_6810 <= 1'h0;
      p11_uge_6888 <= 1'h0;
      p11_uge_6966 <= 1'h0;
      p11_uge_7044 <= 1'h0;
      p11_uge_7122 <= 1'h0;
      p11_uge_7200 <= 1'h0;
      p11_uge_7278 <= 1'h0;
      p11_uge_7356 <= 1'h0;
      p11_uge_7434 <= 1'h0;
      p11_r__22 <= 32'h0000_0000;
      p11_bit_slice_6555 <= 1'h0;
      p11_bit_slice_6556 <= 1'h0;
      p11_bit_slice_6557 <= 1'h0;
      p11_bit_slice_6558 <= 1'h0;
      p11_bit_slice_6559 <= 1'h0;
      p11_bit_slice_6560 <= 1'h0;
      p11_bit_slice_6561 <= 1'h0;
      p11_bit_slice_6562 <= 1'h0;
      p11_bit_slice_6563 <= 1'h0;
      p11_bit_slice_6564 <= 1'h0;
      p11_bit_slice_6565 <= 1'h0;
      p11_bit_slice_6566 <= 1'h0;
      p11_bit_slice_6567 <= 1'h0;
      p11_bit_slice_6568 <= 1'h0;
      p11_bit_slice_6569 <= 1'h0;
      p11_bit_slice_6570 <= 1'h0;
      p11_bit_slice_6571 <= 1'h0;
      p11_bit_slice_6572 <= 1'h0;
      p11_bit_slice_6573 <= 1'h0;
      p11_bit_slice_6574 <= 1'h0;
      p11_bit_slice_6575 <= 1'h0;
      p12_b <= 32'h0000_0000;
      p12_uge_6652 <= 1'h0;
      p12_bivisor__1 <= 33'h0_0000_0000;
      p12_uge_6732 <= 1'h0;
      p12_uge_6810 <= 1'h0;
      p12_uge_6888 <= 1'h0;
      p12_uge_6966 <= 1'h0;
      p12_uge_7044 <= 1'h0;
      p12_uge_7122 <= 1'h0;
      p12_uge_7200 <= 1'h0;
      p12_uge_7278 <= 1'h0;
      p12_uge_7356 <= 1'h0;
      p12_uge_7434 <= 1'h0;
      p12_uge_7512 <= 1'h0;
      p12_r__24 <= 32'h0000_0000;
      p12_bit_slice_6556 <= 1'h0;
      p12_bit_slice_6557 <= 1'h0;
      p12_bit_slice_6558 <= 1'h0;
      p12_bit_slice_6559 <= 1'h0;
      p12_bit_slice_6560 <= 1'h0;
      p12_bit_slice_6561 <= 1'h0;
      p12_bit_slice_6562 <= 1'h0;
      p12_bit_slice_6563 <= 1'h0;
      p12_bit_slice_6564 <= 1'h0;
      p12_bit_slice_6565 <= 1'h0;
      p12_bit_slice_6566 <= 1'h0;
      p12_bit_slice_6567 <= 1'h0;
      p12_bit_slice_6568 <= 1'h0;
      p12_bit_slice_6569 <= 1'h0;
      p12_bit_slice_6570 <= 1'h0;
      p12_bit_slice_6571 <= 1'h0;
      p12_bit_slice_6572 <= 1'h0;
      p12_bit_slice_6573 <= 1'h0;
      p12_bit_slice_6574 <= 1'h0;
      p12_bit_slice_6575 <= 1'h0;
      p13_b <= 32'h0000_0000;
      p13_uge_6652 <= 1'h0;
      p13_bivisor__1 <= 33'h0_0000_0000;
      p13_uge_6732 <= 1'h0;
      p13_uge_6810 <= 1'h0;
      p13_uge_6888 <= 1'h0;
      p13_uge_6966 <= 1'h0;
      p13_uge_7044 <= 1'h0;
      p13_uge_7122 <= 1'h0;
      p13_uge_7200 <= 1'h0;
      p13_uge_7278 <= 1'h0;
      p13_uge_7356 <= 1'h0;
      p13_uge_7434 <= 1'h0;
      p13_uge_7512 <= 1'h0;
      p13_uge_7590 <= 1'h0;
      p13_r__26 <= 32'h0000_0000;
      p13_bit_slice_6557 <= 1'h0;
      p13_bit_slice_6558 <= 1'h0;
      p13_bit_slice_6559 <= 1'h0;
      p13_bit_slice_6560 <= 1'h0;
      p13_bit_slice_6561 <= 1'h0;
      p13_bit_slice_6562 <= 1'h0;
      p13_bit_slice_6563 <= 1'h0;
      p13_bit_slice_6564 <= 1'h0;
      p13_bit_slice_6565 <= 1'h0;
      p13_bit_slice_6566 <= 1'h0;
      p13_bit_slice_6567 <= 1'h0;
      p13_bit_slice_6568 <= 1'h0;
      p13_bit_slice_6569 <= 1'h0;
      p13_bit_slice_6570 <= 1'h0;
      p13_bit_slice_6571 <= 1'h0;
      p13_bit_slice_6572 <= 1'h0;
      p13_bit_slice_6573 <= 1'h0;
      p13_bit_slice_6574 <= 1'h0;
      p13_bit_slice_6575 <= 1'h0;
      p14_b <= 32'h0000_0000;
      p14_uge_6652 <= 1'h0;
      p14_bivisor__1 <= 33'h0_0000_0000;
      p14_uge_6732 <= 1'h0;
      p14_uge_6810 <= 1'h0;
      p14_uge_6888 <= 1'h0;
      p14_uge_6966 <= 1'h0;
      p14_uge_7044 <= 1'h0;
      p14_uge_7122 <= 1'h0;
      p14_uge_7200 <= 1'h0;
      p14_uge_7278 <= 1'h0;
      p14_uge_7356 <= 1'h0;
      p14_uge_7434 <= 1'h0;
      p14_uge_7512 <= 1'h0;
      p14_uge_7590 <= 1'h0;
      p14_uge_7668 <= 1'h0;
      p14_r__28 <= 32'h0000_0000;
      p14_bit_slice_6558 <= 1'h0;
      p14_bit_slice_6559 <= 1'h0;
      p14_bit_slice_6560 <= 1'h0;
      p14_bit_slice_6561 <= 1'h0;
      p14_bit_slice_6562 <= 1'h0;
      p14_bit_slice_6563 <= 1'h0;
      p14_bit_slice_6564 <= 1'h0;
      p14_bit_slice_6565 <= 1'h0;
      p14_bit_slice_6566 <= 1'h0;
      p14_bit_slice_6567 <= 1'h0;
      p14_bit_slice_6568 <= 1'h0;
      p14_bit_slice_6569 <= 1'h0;
      p14_bit_slice_6570 <= 1'h0;
      p14_bit_slice_6571 <= 1'h0;
      p14_bit_slice_6572 <= 1'h0;
      p14_bit_slice_6573 <= 1'h0;
      p14_bit_slice_6574 <= 1'h0;
      p14_bit_slice_6575 <= 1'h0;
      p15_b <= 32'h0000_0000;
      p15_uge_6652 <= 1'h0;
      p15_bivisor__1 <= 33'h0_0000_0000;
      p15_uge_6732 <= 1'h0;
      p15_uge_6810 <= 1'h0;
      p15_uge_6888 <= 1'h0;
      p15_uge_6966 <= 1'h0;
      p15_uge_7044 <= 1'h0;
      p15_uge_7122 <= 1'h0;
      p15_uge_7200 <= 1'h0;
      p15_uge_7278 <= 1'h0;
      p15_uge_7356 <= 1'h0;
      p15_uge_7434 <= 1'h0;
      p15_uge_7512 <= 1'h0;
      p15_uge_7590 <= 1'h0;
      p15_uge_7668 <= 1'h0;
      p15_uge_7746 <= 1'h0;
      p15_r__30 <= 32'h0000_0000;
      p15_bit_slice_6559 <= 1'h0;
      p15_bit_slice_6560 <= 1'h0;
      p15_bit_slice_6561 <= 1'h0;
      p15_bit_slice_6562 <= 1'h0;
      p15_bit_slice_6563 <= 1'h0;
      p15_bit_slice_6564 <= 1'h0;
      p15_bit_slice_6565 <= 1'h0;
      p15_bit_slice_6566 <= 1'h0;
      p15_bit_slice_6567 <= 1'h0;
      p15_bit_slice_6568 <= 1'h0;
      p15_bit_slice_6569 <= 1'h0;
      p15_bit_slice_6570 <= 1'h0;
      p15_bit_slice_6571 <= 1'h0;
      p15_bit_slice_6572 <= 1'h0;
      p15_bit_slice_6573 <= 1'h0;
      p15_bit_slice_6574 <= 1'h0;
      p15_bit_slice_6575 <= 1'h0;
      p16_b <= 32'h0000_0000;
      p16_uge_6652 <= 1'h0;
      p16_bivisor__1 <= 33'h0_0000_0000;
      p16_uge_6732 <= 1'h0;
      p16_uge_6810 <= 1'h0;
      p16_uge_6888 <= 1'h0;
      p16_uge_6966 <= 1'h0;
      p16_uge_7044 <= 1'h0;
      p16_uge_7122 <= 1'h0;
      p16_uge_7200 <= 1'h0;
      p16_uge_7278 <= 1'h0;
      p16_uge_7356 <= 1'h0;
      p16_uge_7434 <= 1'h0;
      p16_uge_7512 <= 1'h0;
      p16_uge_7590 <= 1'h0;
      p16_uge_7668 <= 1'h0;
      p16_uge_7746 <= 1'h0;
      p16_uge_7824 <= 1'h0;
      p16_r__32 <= 32'h0000_0000;
      p16_bit_slice_6560 <= 1'h0;
      p16_bit_slice_6561 <= 1'h0;
      p16_bit_slice_6562 <= 1'h0;
      p16_bit_slice_6563 <= 1'h0;
      p16_bit_slice_6564 <= 1'h0;
      p16_bit_slice_6565 <= 1'h0;
      p16_bit_slice_6566 <= 1'h0;
      p16_bit_slice_6567 <= 1'h0;
      p16_bit_slice_6568 <= 1'h0;
      p16_bit_slice_6569 <= 1'h0;
      p16_bit_slice_6570 <= 1'h0;
      p16_bit_slice_6571 <= 1'h0;
      p16_bit_slice_6572 <= 1'h0;
      p16_bit_slice_6573 <= 1'h0;
      p16_bit_slice_6574 <= 1'h0;
      p16_bit_slice_6575 <= 1'h0;
      p17_b <= 32'h0000_0000;
      p17_uge_6652 <= 1'h0;
      p17_bivisor__1 <= 33'h0_0000_0000;
      p17_uge_6732 <= 1'h0;
      p17_uge_6810 <= 1'h0;
      p17_uge_6888 <= 1'h0;
      p17_uge_6966 <= 1'h0;
      p17_uge_7044 <= 1'h0;
      p17_uge_7122 <= 1'h0;
      p17_uge_7200 <= 1'h0;
      p17_uge_7278 <= 1'h0;
      p17_uge_7356 <= 1'h0;
      p17_uge_7434 <= 1'h0;
      p17_uge_7512 <= 1'h0;
      p17_uge_7590 <= 1'h0;
      p17_uge_7668 <= 1'h0;
      p17_uge_7746 <= 1'h0;
      p17_uge_7824 <= 1'h0;
      p17_uge_7902 <= 1'h0;
      p17_r__34 <= 32'h0000_0000;
      p17_bit_slice_6561 <= 1'h0;
      p17_bit_slice_6562 <= 1'h0;
      p17_bit_slice_6563 <= 1'h0;
      p17_bit_slice_6564 <= 1'h0;
      p17_bit_slice_6565 <= 1'h0;
      p17_bit_slice_6566 <= 1'h0;
      p17_bit_slice_6567 <= 1'h0;
      p17_bit_slice_6568 <= 1'h0;
      p17_bit_slice_6569 <= 1'h0;
      p17_bit_slice_6570 <= 1'h0;
      p17_bit_slice_6571 <= 1'h0;
      p17_bit_slice_6572 <= 1'h0;
      p17_bit_slice_6573 <= 1'h0;
      p17_bit_slice_6574 <= 1'h0;
      p17_bit_slice_6575 <= 1'h0;
      p18_b <= 32'h0000_0000;
      p18_uge_6652 <= 1'h0;
      p18_bivisor__1 <= 33'h0_0000_0000;
      p18_uge_6732 <= 1'h0;
      p18_uge_6810 <= 1'h0;
      p18_uge_6888 <= 1'h0;
      p18_uge_6966 <= 1'h0;
      p18_uge_7044 <= 1'h0;
      p18_uge_7122 <= 1'h0;
      p18_uge_7200 <= 1'h0;
      p18_uge_7278 <= 1'h0;
      p18_uge_7356 <= 1'h0;
      p18_uge_7434 <= 1'h0;
      p18_uge_7512 <= 1'h0;
      p18_uge_7590 <= 1'h0;
      p18_uge_7668 <= 1'h0;
      p18_uge_7746 <= 1'h0;
      p18_uge_7824 <= 1'h0;
      p18_uge_7902 <= 1'h0;
      p18_uge_7980 <= 1'h0;
      p18_r__36 <= 32'h0000_0000;
      p18_bit_slice_6562 <= 1'h0;
      p18_bit_slice_6563 <= 1'h0;
      p18_bit_slice_6564 <= 1'h0;
      p18_bit_slice_6565 <= 1'h0;
      p18_bit_slice_6566 <= 1'h0;
      p18_bit_slice_6567 <= 1'h0;
      p18_bit_slice_6568 <= 1'h0;
      p18_bit_slice_6569 <= 1'h0;
      p18_bit_slice_6570 <= 1'h0;
      p18_bit_slice_6571 <= 1'h0;
      p18_bit_slice_6572 <= 1'h0;
      p18_bit_slice_6573 <= 1'h0;
      p18_bit_slice_6574 <= 1'h0;
      p18_bit_slice_6575 <= 1'h0;
      p19_b <= 32'h0000_0000;
      p19_uge_6652 <= 1'h0;
      p19_bivisor__1 <= 33'h0_0000_0000;
      p19_uge_6732 <= 1'h0;
      p19_uge_6810 <= 1'h0;
      p19_uge_6888 <= 1'h0;
      p19_uge_6966 <= 1'h0;
      p19_uge_7044 <= 1'h0;
      p19_uge_7122 <= 1'h0;
      p19_uge_7200 <= 1'h0;
      p19_uge_7278 <= 1'h0;
      p19_uge_7356 <= 1'h0;
      p19_uge_7434 <= 1'h0;
      p19_uge_7512 <= 1'h0;
      p19_uge_7590 <= 1'h0;
      p19_uge_7668 <= 1'h0;
      p19_uge_7746 <= 1'h0;
      p19_uge_7824 <= 1'h0;
      p19_uge_7902 <= 1'h0;
      p19_uge_7980 <= 1'h0;
      p19_uge_8058 <= 1'h0;
      p19_r__38 <= 32'h0000_0000;
      p19_bit_slice_6563 <= 1'h0;
      p19_bit_slice_6564 <= 1'h0;
      p19_bit_slice_6565 <= 1'h0;
      p19_bit_slice_6566 <= 1'h0;
      p19_bit_slice_6567 <= 1'h0;
      p19_bit_slice_6568 <= 1'h0;
      p19_bit_slice_6569 <= 1'h0;
      p19_bit_slice_6570 <= 1'h0;
      p19_bit_slice_6571 <= 1'h0;
      p19_bit_slice_6572 <= 1'h0;
      p19_bit_slice_6573 <= 1'h0;
      p19_bit_slice_6574 <= 1'h0;
      p19_bit_slice_6575 <= 1'h0;
      p20_b <= 32'h0000_0000;
      p20_uge_6652 <= 1'h0;
      p20_bivisor__1 <= 33'h0_0000_0000;
      p20_uge_6732 <= 1'h0;
      p20_uge_6810 <= 1'h0;
      p20_uge_6888 <= 1'h0;
      p20_uge_6966 <= 1'h0;
      p20_uge_7044 <= 1'h0;
      p20_uge_7122 <= 1'h0;
      p20_uge_7200 <= 1'h0;
      p20_uge_7278 <= 1'h0;
      p20_uge_7356 <= 1'h0;
      p20_uge_7434 <= 1'h0;
      p20_uge_7512 <= 1'h0;
      p20_uge_7590 <= 1'h0;
      p20_uge_7668 <= 1'h0;
      p20_uge_7746 <= 1'h0;
      p20_uge_7824 <= 1'h0;
      p20_uge_7902 <= 1'h0;
      p20_uge_7980 <= 1'h0;
      p20_uge_8058 <= 1'h0;
      p20_uge_8136 <= 1'h0;
      p20_r__40 <= 32'h0000_0000;
      p20_bit_slice_6564 <= 1'h0;
      p20_bit_slice_6565 <= 1'h0;
      p20_bit_slice_6566 <= 1'h0;
      p20_bit_slice_6567 <= 1'h0;
      p20_bit_slice_6568 <= 1'h0;
      p20_bit_slice_6569 <= 1'h0;
      p20_bit_slice_6570 <= 1'h0;
      p20_bit_slice_6571 <= 1'h0;
      p20_bit_slice_6572 <= 1'h0;
      p20_bit_slice_6573 <= 1'h0;
      p20_bit_slice_6574 <= 1'h0;
      p20_bit_slice_6575 <= 1'h0;
      p21_b <= 32'h0000_0000;
      p21_uge_6652 <= 1'h0;
      p21_bivisor__1 <= 33'h0_0000_0000;
      p21_uge_6732 <= 1'h0;
      p21_uge_6810 <= 1'h0;
      p21_uge_6888 <= 1'h0;
      p21_uge_6966 <= 1'h0;
      p21_uge_7044 <= 1'h0;
      p21_uge_7122 <= 1'h0;
      p21_uge_7200 <= 1'h0;
      p21_uge_7278 <= 1'h0;
      p21_uge_7356 <= 1'h0;
      p21_uge_7434 <= 1'h0;
      p21_uge_7512 <= 1'h0;
      p21_uge_7590 <= 1'h0;
      p21_uge_7668 <= 1'h0;
      p21_uge_7746 <= 1'h0;
      p21_uge_7824 <= 1'h0;
      p21_uge_7902 <= 1'h0;
      p21_uge_7980 <= 1'h0;
      p21_uge_8058 <= 1'h0;
      p21_uge_8136 <= 1'h0;
      p21_uge_8214 <= 1'h0;
      p21_r__42 <= 32'h0000_0000;
      p21_bit_slice_6565 <= 1'h0;
      p21_bit_slice_6566 <= 1'h0;
      p21_bit_slice_6567 <= 1'h0;
      p21_bit_slice_6568 <= 1'h0;
      p21_bit_slice_6569 <= 1'h0;
      p21_bit_slice_6570 <= 1'h0;
      p21_bit_slice_6571 <= 1'h0;
      p21_bit_slice_6572 <= 1'h0;
      p21_bit_slice_6573 <= 1'h0;
      p21_bit_slice_6574 <= 1'h0;
      p21_bit_slice_6575 <= 1'h0;
      p22_b <= 32'h0000_0000;
      p22_uge_6652 <= 1'h0;
      p22_bivisor__1 <= 33'h0_0000_0000;
      p22_uge_6732 <= 1'h0;
      p22_uge_6810 <= 1'h0;
      p22_uge_6888 <= 1'h0;
      p22_uge_6966 <= 1'h0;
      p22_uge_7044 <= 1'h0;
      p22_uge_7122 <= 1'h0;
      p22_uge_7200 <= 1'h0;
      p22_uge_7278 <= 1'h0;
      p22_uge_7356 <= 1'h0;
      p22_uge_7434 <= 1'h0;
      p22_uge_7512 <= 1'h0;
      p22_uge_7590 <= 1'h0;
      p22_uge_7668 <= 1'h0;
      p22_uge_7746 <= 1'h0;
      p22_uge_7824 <= 1'h0;
      p22_uge_7902 <= 1'h0;
      p22_uge_7980 <= 1'h0;
      p22_uge_8058 <= 1'h0;
      p22_uge_8136 <= 1'h0;
      p22_uge_8214 <= 1'h0;
      p22_uge_8292 <= 1'h0;
      p22_r__44 <= 32'h0000_0000;
      p22_bit_slice_6566 <= 1'h0;
      p22_bit_slice_6567 <= 1'h0;
      p22_bit_slice_6568 <= 1'h0;
      p22_bit_slice_6569 <= 1'h0;
      p22_bit_slice_6570 <= 1'h0;
      p22_bit_slice_6571 <= 1'h0;
      p22_bit_slice_6572 <= 1'h0;
      p22_bit_slice_6573 <= 1'h0;
      p22_bit_slice_6574 <= 1'h0;
      p22_bit_slice_6575 <= 1'h0;
      p23_b <= 32'h0000_0000;
      p23_uge_6652 <= 1'h0;
      p23_bivisor__1 <= 33'h0_0000_0000;
      p23_uge_6732 <= 1'h0;
      p23_uge_6810 <= 1'h0;
      p23_uge_6888 <= 1'h0;
      p23_uge_6966 <= 1'h0;
      p23_uge_7044 <= 1'h0;
      p23_uge_7122 <= 1'h0;
      p23_uge_7200 <= 1'h0;
      p23_uge_7278 <= 1'h0;
      p23_uge_7356 <= 1'h0;
      p23_uge_7434 <= 1'h0;
      p23_uge_7512 <= 1'h0;
      p23_uge_7590 <= 1'h0;
      p23_uge_7668 <= 1'h0;
      p23_uge_7746 <= 1'h0;
      p23_uge_7824 <= 1'h0;
      p23_uge_7902 <= 1'h0;
      p23_uge_7980 <= 1'h0;
      p23_uge_8058 <= 1'h0;
      p23_uge_8136 <= 1'h0;
      p23_uge_8214 <= 1'h0;
      p23_uge_8292 <= 1'h0;
      p23_uge_8370 <= 1'h0;
      p23_r__46 <= 32'h0000_0000;
      p23_bit_slice_6567 <= 1'h0;
      p23_bit_slice_6568 <= 1'h0;
      p23_bit_slice_6569 <= 1'h0;
      p23_bit_slice_6570 <= 1'h0;
      p23_bit_slice_6571 <= 1'h0;
      p23_bit_slice_6572 <= 1'h0;
      p23_bit_slice_6573 <= 1'h0;
      p23_bit_slice_6574 <= 1'h0;
      p23_bit_slice_6575 <= 1'h0;
      p24_b <= 32'h0000_0000;
      p24_uge_6652 <= 1'h0;
      p24_bivisor__1 <= 33'h0_0000_0000;
      p24_uge_6732 <= 1'h0;
      p24_uge_6810 <= 1'h0;
      p24_uge_6888 <= 1'h0;
      p24_uge_6966 <= 1'h0;
      p24_uge_7044 <= 1'h0;
      p24_uge_7122 <= 1'h0;
      p24_uge_7200 <= 1'h0;
      p24_uge_7278 <= 1'h0;
      p24_uge_7356 <= 1'h0;
      p24_uge_7434 <= 1'h0;
      p24_uge_7512 <= 1'h0;
      p24_uge_7590 <= 1'h0;
      p24_uge_7668 <= 1'h0;
      p24_uge_7746 <= 1'h0;
      p24_uge_7824 <= 1'h0;
      p24_uge_7902 <= 1'h0;
      p24_uge_7980 <= 1'h0;
      p24_uge_8058 <= 1'h0;
      p24_uge_8136 <= 1'h0;
      p24_uge_8214 <= 1'h0;
      p24_uge_8292 <= 1'h0;
      p24_uge_8370 <= 1'h0;
      p24_uge_8448 <= 1'h0;
      p24_r__48 <= 32'h0000_0000;
      p24_bit_slice_6568 <= 1'h0;
      p24_bit_slice_6569 <= 1'h0;
      p24_bit_slice_6570 <= 1'h0;
      p24_bit_slice_6571 <= 1'h0;
      p24_bit_slice_6572 <= 1'h0;
      p24_bit_slice_6573 <= 1'h0;
      p24_bit_slice_6574 <= 1'h0;
      p24_bit_slice_6575 <= 1'h0;
      p25_b <= 32'h0000_0000;
      p25_uge_6652 <= 1'h0;
      p25_bivisor__1 <= 33'h0_0000_0000;
      p25_uge_6732 <= 1'h0;
      p25_uge_6810 <= 1'h0;
      p25_uge_6888 <= 1'h0;
      p25_uge_6966 <= 1'h0;
      p25_uge_7044 <= 1'h0;
      p25_uge_7122 <= 1'h0;
      p25_uge_7200 <= 1'h0;
      p25_uge_7278 <= 1'h0;
      p25_uge_7356 <= 1'h0;
      p25_uge_7434 <= 1'h0;
      p25_uge_7512 <= 1'h0;
      p25_uge_7590 <= 1'h0;
      p25_uge_7668 <= 1'h0;
      p25_uge_7746 <= 1'h0;
      p25_uge_7824 <= 1'h0;
      p25_uge_7902 <= 1'h0;
      p25_uge_7980 <= 1'h0;
      p25_uge_8058 <= 1'h0;
      p25_uge_8136 <= 1'h0;
      p25_uge_8214 <= 1'h0;
      p25_uge_8292 <= 1'h0;
      p25_uge_8370 <= 1'h0;
      p25_uge_8448 <= 1'h0;
      p25_uge_8526 <= 1'h0;
      p25_r__50 <= 32'h0000_0000;
      p25_bit_slice_6569 <= 1'h0;
      p25_bit_slice_6570 <= 1'h0;
      p25_bit_slice_6571 <= 1'h0;
      p25_bit_slice_6572 <= 1'h0;
      p25_bit_slice_6573 <= 1'h0;
      p25_bit_slice_6574 <= 1'h0;
      p25_bit_slice_6575 <= 1'h0;
      p26_b <= 32'h0000_0000;
      p26_uge_6652 <= 1'h0;
      p26_bivisor__1 <= 33'h0_0000_0000;
      p26_uge_6732 <= 1'h0;
      p26_uge_6810 <= 1'h0;
      p26_uge_6888 <= 1'h0;
      p26_uge_6966 <= 1'h0;
      p26_uge_7044 <= 1'h0;
      p26_uge_7122 <= 1'h0;
      p26_uge_7200 <= 1'h0;
      p26_uge_7278 <= 1'h0;
      p26_uge_7356 <= 1'h0;
      p26_uge_7434 <= 1'h0;
      p26_uge_7512 <= 1'h0;
      p26_uge_7590 <= 1'h0;
      p26_uge_7668 <= 1'h0;
      p26_uge_7746 <= 1'h0;
      p26_uge_7824 <= 1'h0;
      p26_uge_7902 <= 1'h0;
      p26_uge_7980 <= 1'h0;
      p26_uge_8058 <= 1'h0;
      p26_uge_8136 <= 1'h0;
      p26_uge_8214 <= 1'h0;
      p26_uge_8292 <= 1'h0;
      p26_uge_8370 <= 1'h0;
      p26_uge_8448 <= 1'h0;
      p26_uge_8526 <= 1'h0;
      p26_uge_8604 <= 1'h0;
      p26_r__52 <= 32'h0000_0000;
      p26_bit_slice_6570 <= 1'h0;
      p26_bit_slice_6571 <= 1'h0;
      p26_bit_slice_6572 <= 1'h0;
      p26_bit_slice_6573 <= 1'h0;
      p26_bit_slice_6574 <= 1'h0;
      p26_bit_slice_6575 <= 1'h0;
      p27_b <= 32'h0000_0000;
      p27_uge_6652 <= 1'h0;
      p27_bivisor__1 <= 33'h0_0000_0000;
      p27_uge_6732 <= 1'h0;
      p27_uge_6810 <= 1'h0;
      p27_uge_6888 <= 1'h0;
      p27_uge_6966 <= 1'h0;
      p27_uge_7044 <= 1'h0;
      p27_uge_7122 <= 1'h0;
      p27_uge_7200 <= 1'h0;
      p27_uge_7278 <= 1'h0;
      p27_uge_7356 <= 1'h0;
      p27_uge_7434 <= 1'h0;
      p27_uge_7512 <= 1'h0;
      p27_uge_7590 <= 1'h0;
      p27_uge_7668 <= 1'h0;
      p27_uge_7746 <= 1'h0;
      p27_uge_7824 <= 1'h0;
      p27_uge_7902 <= 1'h0;
      p27_uge_7980 <= 1'h0;
      p27_uge_8058 <= 1'h0;
      p27_uge_8136 <= 1'h0;
      p27_uge_8214 <= 1'h0;
      p27_uge_8292 <= 1'h0;
      p27_uge_8370 <= 1'h0;
      p27_uge_8448 <= 1'h0;
      p27_uge_8526 <= 1'h0;
      p27_uge_8604 <= 1'h0;
      p27_uge_8682 <= 1'h0;
      p27_r__54 <= 32'h0000_0000;
      p27_bit_slice_6571 <= 1'h0;
      p27_bit_slice_6572 <= 1'h0;
      p27_bit_slice_6573 <= 1'h0;
      p27_bit_slice_6574 <= 1'h0;
      p27_bit_slice_6575 <= 1'h0;
      p28_b <= 32'h0000_0000;
      p28_uge_6652 <= 1'h0;
      p28_bivisor__1 <= 33'h0_0000_0000;
      p28_uge_6732 <= 1'h0;
      p28_uge_6810 <= 1'h0;
      p28_uge_6888 <= 1'h0;
      p28_uge_6966 <= 1'h0;
      p28_uge_7044 <= 1'h0;
      p28_uge_7122 <= 1'h0;
      p28_uge_7200 <= 1'h0;
      p28_uge_7278 <= 1'h0;
      p28_uge_7356 <= 1'h0;
      p28_uge_7434 <= 1'h0;
      p28_uge_7512 <= 1'h0;
      p28_uge_7590 <= 1'h0;
      p28_uge_7668 <= 1'h0;
      p28_uge_7746 <= 1'h0;
      p28_uge_7824 <= 1'h0;
      p28_uge_7902 <= 1'h0;
      p28_uge_7980 <= 1'h0;
      p28_uge_8058 <= 1'h0;
      p28_uge_8136 <= 1'h0;
      p28_uge_8214 <= 1'h0;
      p28_uge_8292 <= 1'h0;
      p28_uge_8370 <= 1'h0;
      p28_uge_8448 <= 1'h0;
      p28_uge_8526 <= 1'h0;
      p28_uge_8604 <= 1'h0;
      p28_uge_8682 <= 1'h0;
      p28_uge_8760 <= 1'h0;
      p28_r__56 <= 32'h0000_0000;
      p28_bit_slice_6572 <= 1'h0;
      p28_bit_slice_6573 <= 1'h0;
      p28_bit_slice_6574 <= 1'h0;
      p28_bit_slice_6575 <= 1'h0;
      p29_b <= 32'h0000_0000;
      p29_uge_6652 <= 1'h0;
      p29_bivisor__1 <= 33'h0_0000_0000;
      p29_uge_6732 <= 1'h0;
      p29_uge_6810 <= 1'h0;
      p29_uge_6888 <= 1'h0;
      p29_uge_6966 <= 1'h0;
      p29_uge_7044 <= 1'h0;
      p29_uge_7122 <= 1'h0;
      p29_uge_7200 <= 1'h0;
      p29_uge_7278 <= 1'h0;
      p29_uge_7356 <= 1'h0;
      p29_uge_7434 <= 1'h0;
      p29_uge_7512 <= 1'h0;
      p29_uge_7590 <= 1'h0;
      p29_uge_7668 <= 1'h0;
      p29_uge_7746 <= 1'h0;
      p29_uge_7824 <= 1'h0;
      p29_uge_7902 <= 1'h0;
      p29_uge_7980 <= 1'h0;
      p29_uge_8058 <= 1'h0;
      p29_uge_8136 <= 1'h0;
      p29_uge_8214 <= 1'h0;
      p29_uge_8292 <= 1'h0;
      p29_uge_8370 <= 1'h0;
      p29_uge_8448 <= 1'h0;
      p29_uge_8526 <= 1'h0;
      p29_uge_8604 <= 1'h0;
      p29_uge_8682 <= 1'h0;
      p29_uge_8760 <= 1'h0;
      p29_uge_8838 <= 1'h0;
      p29_r__58 <= 32'h0000_0000;
      p29_bit_slice_6573 <= 1'h0;
      p29_bit_slice_6574 <= 1'h0;
      p29_bit_slice_6575 <= 1'h0;
      p30_b <= 32'h0000_0000;
      p30_uge_6652 <= 1'h0;
      p30_bivisor__1 <= 33'h0_0000_0000;
      p30_uge_6732 <= 1'h0;
      p30_uge_6810 <= 1'h0;
      p30_uge_6888 <= 1'h0;
      p30_uge_6966 <= 1'h0;
      p30_uge_7044 <= 1'h0;
      p30_uge_7122 <= 1'h0;
      p30_uge_7200 <= 1'h0;
      p30_uge_7278 <= 1'h0;
      p30_uge_7356 <= 1'h0;
      p30_uge_7434 <= 1'h0;
      p30_uge_7512 <= 1'h0;
      p30_uge_7590 <= 1'h0;
      p30_uge_7668 <= 1'h0;
      p30_uge_7746 <= 1'h0;
      p30_uge_7824 <= 1'h0;
      p30_uge_7902 <= 1'h0;
      p30_uge_7980 <= 1'h0;
      p30_uge_8058 <= 1'h0;
      p30_uge_8136 <= 1'h0;
      p30_uge_8214 <= 1'h0;
      p30_uge_8292 <= 1'h0;
      p30_uge_8370 <= 1'h0;
      p30_uge_8448 <= 1'h0;
      p30_uge_8526 <= 1'h0;
      p30_uge_8604 <= 1'h0;
      p30_uge_8682 <= 1'h0;
      p30_uge_8760 <= 1'h0;
      p30_uge_8838 <= 1'h0;
      p30_uge_8916 <= 1'h0;
      p30_r__60 <= 32'h0000_0000;
      p30_bit_slice_6574 <= 1'h0;
      p30_bit_slice_6575 <= 1'h0;
      p31_uge_6652 <= 1'h0;
      p31_bivisor__1 <= 33'h0_0000_0000;
      p31_uge_6732 <= 1'h0;
      p31_uge_6810 <= 1'h0;
      p31_uge_6888 <= 1'h0;
      p31_uge_6966 <= 1'h0;
      p31_uge_7044 <= 1'h0;
      p31_uge_7122 <= 1'h0;
      p31_uge_7200 <= 1'h0;
      p31_uge_7278 <= 1'h0;
      p31_uge_7356 <= 1'h0;
      p31_uge_7434 <= 1'h0;
      p31_uge_7512 <= 1'h0;
      p31_uge_7590 <= 1'h0;
      p31_uge_7668 <= 1'h0;
      p31_uge_7746 <= 1'h0;
      p31_uge_7824 <= 1'h0;
      p31_uge_7902 <= 1'h0;
      p31_uge_7980 <= 1'h0;
      p31_uge_8058 <= 1'h0;
      p31_uge_8136 <= 1'h0;
      p31_uge_8214 <= 1'h0;
      p31_uge_8292 <= 1'h0;
      p31_uge_8370 <= 1'h0;
      p31_uge_8448 <= 1'h0;
      p31_uge_8526 <= 1'h0;
      p31_uge_8604 <= 1'h0;
      p31_uge_8682 <= 1'h0;
      p31_uge_8760 <= 1'h0;
      p31_uge_8838 <= 1'h0;
      p31_uge_8916 <= 1'h0;
      p31_uge_8994 <= 1'h0;
      p31_r__62 <= 32'h0000_0000;
      p31_bit_slice_6575 <= 1'h0;
      p0_valid <= 1'h0;
      p1_valid <= 1'h0;
      p2_valid <= 1'h0;
      p3_valid <= 1'h0;
      p4_valid <= 1'h0;
      p5_valid <= 1'h0;
      p6_valid <= 1'h0;
      p7_valid <= 1'h0;
      p8_valid <= 1'h0;
      p9_valid <= 1'h0;
      p10_valid <= 1'h0;
      p11_valid <= 1'h0;
      p12_valid <= 1'h0;
      p13_valid <= 1'h0;
      p14_valid <= 1'h0;
      p15_valid <= 1'h0;
      p16_valid <= 1'h0;
      p17_valid <= 1'h0;
      p18_valid <= 1'h0;
      p19_valid <= 1'h0;
      p20_valid <= 1'h0;
      p21_valid <= 1'h0;
      p22_valid <= 1'h0;
      p23_valid <= 1'h0;
      p24_valid <= 1'h0;
      p25_valid <= 1'h0;
      p26_valid <= 1'h0;
      p27_valid <= 1'h0;
      p28_valid <= 1'h0;
      p29_valid <= 1'h0;
      p30_valid <= 1'h0;
      p31_valid <= 1'h0;
      p32_valid <= 1'h0;
      p33_valid <= 1'h0;
      p34_valid <= 1'h0;
      __xls_float_ips__result_reg <= 32'h0000_0000;
      __xls_float_ips__result_valid_reg <= 1'h0;
    end else begin
      p0_bit_slice_6544 <= p0_data_enable ? bit_slice_6544 : p0_bit_slice_6544;
      p0_bit_slice_6545 <= p0_data_enable ? bit_slice_6545 : p0_bit_slice_6545;
      p0_bit_slice_6546 <= p0_data_enable ? bit_slice_6546 : p0_bit_slice_6546;
      p0_bit_slice_6547 <= p0_data_enable ? bit_slice_6547 : p0_bit_slice_6547;
      p0_bit_slice_6548 <= p0_data_enable ? bit_slice_6548 : p0_bit_slice_6548;
      p0_bit_slice_6549 <= p0_data_enable ? bit_slice_6549 : p0_bit_slice_6549;
      p0_bit_slice_6550 <= p0_data_enable ? bit_slice_6550 : p0_bit_slice_6550;
      p0_bit_slice_6551 <= p0_data_enable ? bit_slice_6551 : p0_bit_slice_6551;
      p0_bit_slice_6552 <= p0_data_enable ? bit_slice_6552 : p0_bit_slice_6552;
      p0_bit_slice_6553 <= p0_data_enable ? bit_slice_6553 : p0_bit_slice_6553;
      p0_bit_slice_6554 <= p0_data_enable ? bit_slice_6554 : p0_bit_slice_6554;
      p0_bit_slice_6555 <= p0_data_enable ? bit_slice_6555 : p0_bit_slice_6555;
      p0_bit_slice_6556 <= p0_data_enable ? bit_slice_6556 : p0_bit_slice_6556;
      p0_bit_slice_6557 <= p0_data_enable ? bit_slice_6557 : p0_bit_slice_6557;
      p0_bit_slice_6558 <= p0_data_enable ? bit_slice_6558 : p0_bit_slice_6558;
      p0_bit_slice_6559 <= p0_data_enable ? bit_slice_6559 : p0_bit_slice_6559;
      p0_bit_slice_6560 <= p0_data_enable ? bit_slice_6560 : p0_bit_slice_6560;
      p0_bit_slice_6561 <= p0_data_enable ? bit_slice_6561 : p0_bit_slice_6561;
      p0_bit_slice_6562 <= p0_data_enable ? bit_slice_6562 : p0_bit_slice_6562;
      p0_bit_slice_6563 <= p0_data_enable ? bit_slice_6563 : p0_bit_slice_6563;
      p0_bit_slice_6564 <= p0_data_enable ? bit_slice_6564 : p0_bit_slice_6564;
      p0_bit_slice_6565 <= p0_data_enable ? bit_slice_6565 : p0_bit_slice_6565;
      p0_bit_slice_6566 <= p0_data_enable ? bit_slice_6566 : p0_bit_slice_6566;
      p0_bit_slice_6567 <= p0_data_enable ? bit_slice_6567 : p0_bit_slice_6567;
      p0_bit_slice_6568 <= p0_data_enable ? bit_slice_6568 : p0_bit_slice_6568;
      p0_bit_slice_6569 <= p0_data_enable ? bit_slice_6569 : p0_bit_slice_6569;
      p0_bit_slice_6570 <= p0_data_enable ? bit_slice_6570 : p0_bit_slice_6570;
      p0_bit_slice_6571 <= p0_data_enable ? bit_slice_6571 : p0_bit_slice_6571;
      p0_bit_slice_6572 <= p0_data_enable ? bit_slice_6572 : p0_bit_slice_6572;
      p0_bit_slice_6573 <= p0_data_enable ? bit_slice_6573 : p0_bit_slice_6573;
      p0_bit_slice_6574 <= p0_data_enable ? bit_slice_6574 : p0_bit_slice_6574;
      p0_bit_slice_6575 <= p0_data_enable ? bit_slice_6575 : p0_bit_slice_6575;
      p1_b <= p1_data_enable ? xls_float_ips__rhs : p1_b;
      p1_uge_6652 <= p1_data_enable ? uge_6652 : p1_uge_6652;
      p1_r__2 <= p1_data_enable ? r__2 : p1_r__2;
      p1_bit_slice_6545 <= p1_data_enable ? p0_bit_slice_6545 : p1_bit_slice_6545;
      p1_bit_slice_6546 <= p1_data_enable ? p0_bit_slice_6546 : p1_bit_slice_6546;
      p1_bit_slice_6547 <= p1_data_enable ? p0_bit_slice_6547 : p1_bit_slice_6547;
      p1_bit_slice_6548 <= p1_data_enable ? p0_bit_slice_6548 : p1_bit_slice_6548;
      p1_bit_slice_6549 <= p1_data_enable ? p0_bit_slice_6549 : p1_bit_slice_6549;
      p1_bit_slice_6550 <= p1_data_enable ? p0_bit_slice_6550 : p1_bit_slice_6550;
      p1_bit_slice_6551 <= p1_data_enable ? p0_bit_slice_6551 : p1_bit_slice_6551;
      p1_bit_slice_6552 <= p1_data_enable ? p0_bit_slice_6552 : p1_bit_slice_6552;
      p1_bit_slice_6553 <= p1_data_enable ? p0_bit_slice_6553 : p1_bit_slice_6553;
      p1_bit_slice_6554 <= p1_data_enable ? p0_bit_slice_6554 : p1_bit_slice_6554;
      p1_bit_slice_6555 <= p1_data_enable ? p0_bit_slice_6555 : p1_bit_slice_6555;
      p1_bit_slice_6556 <= p1_data_enable ? p0_bit_slice_6556 : p1_bit_slice_6556;
      p1_bit_slice_6557 <= p1_data_enable ? p0_bit_slice_6557 : p1_bit_slice_6557;
      p1_bit_slice_6558 <= p1_data_enable ? p0_bit_slice_6558 : p1_bit_slice_6558;
      p1_bit_slice_6559 <= p1_data_enable ? p0_bit_slice_6559 : p1_bit_slice_6559;
      p1_bit_slice_6560 <= p1_data_enable ? p0_bit_slice_6560 : p1_bit_slice_6560;
      p1_bit_slice_6561 <= p1_data_enable ? p0_bit_slice_6561 : p1_bit_slice_6561;
      p1_bit_slice_6562 <= p1_data_enable ? p0_bit_slice_6562 : p1_bit_slice_6562;
      p1_bit_slice_6563 <= p1_data_enable ? p0_bit_slice_6563 : p1_bit_slice_6563;
      p1_bit_slice_6564 <= p1_data_enable ? p0_bit_slice_6564 : p1_bit_slice_6564;
      p1_bit_slice_6565 <= p1_data_enable ? p0_bit_slice_6565 : p1_bit_slice_6565;
      p1_bit_slice_6566 <= p1_data_enable ? p0_bit_slice_6566 : p1_bit_slice_6566;
      p1_bit_slice_6567 <= p1_data_enable ? p0_bit_slice_6567 : p1_bit_slice_6567;
      p1_bit_slice_6568 <= p1_data_enable ? p0_bit_slice_6568 : p1_bit_slice_6568;
      p1_bit_slice_6569 <= p1_data_enable ? p0_bit_slice_6569 : p1_bit_slice_6569;
      p1_bit_slice_6570 <= p1_data_enable ? p0_bit_slice_6570 : p1_bit_slice_6570;
      p1_bit_slice_6571 <= p1_data_enable ? p0_bit_slice_6571 : p1_bit_slice_6571;
      p1_bit_slice_6572 <= p1_data_enable ? p0_bit_slice_6572 : p1_bit_slice_6572;
      p1_bit_slice_6573 <= p1_data_enable ? p0_bit_slice_6573 : p1_bit_slice_6573;
      p1_bit_slice_6574 <= p1_data_enable ? p0_bit_slice_6574 : p1_bit_slice_6574;
      p1_bit_slice_6575 <= p1_data_enable ? p0_bit_slice_6575 : p1_bit_slice_6575;
      p2_b <= p2_data_enable ? p1_b : p2_b;
      p2_uge_6652 <= p2_data_enable ? p1_uge_6652 : p2_uge_6652;
      p2_bivisor__1 <= p2_data_enable ? bivisor__1 : p2_bivisor__1;
      p2_uge_6732 <= p2_data_enable ? uge_6732 : p2_uge_6732;
      p2_r__4 <= p2_data_enable ? r__4 : p2_r__4;
      p2_bit_slice_6546 <= p2_data_enable ? p1_bit_slice_6546 : p2_bit_slice_6546;
      p2_bit_slice_6547 <= p2_data_enable ? p1_bit_slice_6547 : p2_bit_slice_6547;
      p2_bit_slice_6548 <= p2_data_enable ? p1_bit_slice_6548 : p2_bit_slice_6548;
      p2_bit_slice_6549 <= p2_data_enable ? p1_bit_slice_6549 : p2_bit_slice_6549;
      p2_bit_slice_6550 <= p2_data_enable ? p1_bit_slice_6550 : p2_bit_slice_6550;
      p2_bit_slice_6551 <= p2_data_enable ? p1_bit_slice_6551 : p2_bit_slice_6551;
      p2_bit_slice_6552 <= p2_data_enable ? p1_bit_slice_6552 : p2_bit_slice_6552;
      p2_bit_slice_6553 <= p2_data_enable ? p1_bit_slice_6553 : p2_bit_slice_6553;
      p2_bit_slice_6554 <= p2_data_enable ? p1_bit_slice_6554 : p2_bit_slice_6554;
      p2_bit_slice_6555 <= p2_data_enable ? p1_bit_slice_6555 : p2_bit_slice_6555;
      p2_bit_slice_6556 <= p2_data_enable ? p1_bit_slice_6556 : p2_bit_slice_6556;
      p2_bit_slice_6557 <= p2_data_enable ? p1_bit_slice_6557 : p2_bit_slice_6557;
      p2_bit_slice_6558 <= p2_data_enable ? p1_bit_slice_6558 : p2_bit_slice_6558;
      p2_bit_slice_6559 <= p2_data_enable ? p1_bit_slice_6559 : p2_bit_slice_6559;
      p2_bit_slice_6560 <= p2_data_enable ? p1_bit_slice_6560 : p2_bit_slice_6560;
      p2_bit_slice_6561 <= p2_data_enable ? p1_bit_slice_6561 : p2_bit_slice_6561;
      p2_bit_slice_6562 <= p2_data_enable ? p1_bit_slice_6562 : p2_bit_slice_6562;
      p2_bit_slice_6563 <= p2_data_enable ? p1_bit_slice_6563 : p2_bit_slice_6563;
      p2_bit_slice_6564 <= p2_data_enable ? p1_bit_slice_6564 : p2_bit_slice_6564;
      p2_bit_slice_6565 <= p2_data_enable ? p1_bit_slice_6565 : p2_bit_slice_6565;
      p2_bit_slice_6566 <= p2_data_enable ? p1_bit_slice_6566 : p2_bit_slice_6566;
      p2_bit_slice_6567 <= p2_data_enable ? p1_bit_slice_6567 : p2_bit_slice_6567;
      p2_bit_slice_6568 <= p2_data_enable ? p1_bit_slice_6568 : p2_bit_slice_6568;
      p2_bit_slice_6569 <= p2_data_enable ? p1_bit_slice_6569 : p2_bit_slice_6569;
      p2_bit_slice_6570 <= p2_data_enable ? p1_bit_slice_6570 : p2_bit_slice_6570;
      p2_bit_slice_6571 <= p2_data_enable ? p1_bit_slice_6571 : p2_bit_slice_6571;
      p2_bit_slice_6572 <= p2_data_enable ? p1_bit_slice_6572 : p2_bit_slice_6572;
      p2_bit_slice_6573 <= p2_data_enable ? p1_bit_slice_6573 : p2_bit_slice_6573;
      p2_bit_slice_6574 <= p2_data_enable ? p1_bit_slice_6574 : p2_bit_slice_6574;
      p2_bit_slice_6575 <= p2_data_enable ? p1_bit_slice_6575 : p2_bit_slice_6575;
      p3_b <= p3_data_enable ? p2_b : p3_b;
      p3_uge_6652 <= p3_data_enable ? p2_uge_6652 : p3_uge_6652;
      p3_bivisor__1 <= p3_data_enable ? p2_bivisor__1 : p3_bivisor__1;
      p3_uge_6732 <= p3_data_enable ? p2_uge_6732 : p3_uge_6732;
      p3_uge_6810 <= p3_data_enable ? uge_6810 : p3_uge_6810;
      p3_r__6 <= p3_data_enable ? r__6 : p3_r__6;
      p3_bit_slice_6547 <= p3_data_enable ? p2_bit_slice_6547 : p3_bit_slice_6547;
      p3_bit_slice_6548 <= p3_data_enable ? p2_bit_slice_6548 : p3_bit_slice_6548;
      p3_bit_slice_6549 <= p3_data_enable ? p2_bit_slice_6549 : p3_bit_slice_6549;
      p3_bit_slice_6550 <= p3_data_enable ? p2_bit_slice_6550 : p3_bit_slice_6550;
      p3_bit_slice_6551 <= p3_data_enable ? p2_bit_slice_6551 : p3_bit_slice_6551;
      p3_bit_slice_6552 <= p3_data_enable ? p2_bit_slice_6552 : p3_bit_slice_6552;
      p3_bit_slice_6553 <= p3_data_enable ? p2_bit_slice_6553 : p3_bit_slice_6553;
      p3_bit_slice_6554 <= p3_data_enable ? p2_bit_slice_6554 : p3_bit_slice_6554;
      p3_bit_slice_6555 <= p3_data_enable ? p2_bit_slice_6555 : p3_bit_slice_6555;
      p3_bit_slice_6556 <= p3_data_enable ? p2_bit_slice_6556 : p3_bit_slice_6556;
      p3_bit_slice_6557 <= p3_data_enable ? p2_bit_slice_6557 : p3_bit_slice_6557;
      p3_bit_slice_6558 <= p3_data_enable ? p2_bit_slice_6558 : p3_bit_slice_6558;
      p3_bit_slice_6559 <= p3_data_enable ? p2_bit_slice_6559 : p3_bit_slice_6559;
      p3_bit_slice_6560 <= p3_data_enable ? p2_bit_slice_6560 : p3_bit_slice_6560;
      p3_bit_slice_6561 <= p3_data_enable ? p2_bit_slice_6561 : p3_bit_slice_6561;
      p3_bit_slice_6562 <= p3_data_enable ? p2_bit_slice_6562 : p3_bit_slice_6562;
      p3_bit_slice_6563 <= p3_data_enable ? p2_bit_slice_6563 : p3_bit_slice_6563;
      p3_bit_slice_6564 <= p3_data_enable ? p2_bit_slice_6564 : p3_bit_slice_6564;
      p3_bit_slice_6565 <= p3_data_enable ? p2_bit_slice_6565 : p3_bit_slice_6565;
      p3_bit_slice_6566 <= p3_data_enable ? p2_bit_slice_6566 : p3_bit_slice_6566;
      p3_bit_slice_6567 <= p3_data_enable ? p2_bit_slice_6567 : p3_bit_slice_6567;
      p3_bit_slice_6568 <= p3_data_enable ? p2_bit_slice_6568 : p3_bit_slice_6568;
      p3_bit_slice_6569 <= p3_data_enable ? p2_bit_slice_6569 : p3_bit_slice_6569;
      p3_bit_slice_6570 <= p3_data_enable ? p2_bit_slice_6570 : p3_bit_slice_6570;
      p3_bit_slice_6571 <= p3_data_enable ? p2_bit_slice_6571 : p3_bit_slice_6571;
      p3_bit_slice_6572 <= p3_data_enable ? p2_bit_slice_6572 : p3_bit_slice_6572;
      p3_bit_slice_6573 <= p3_data_enable ? p2_bit_slice_6573 : p3_bit_slice_6573;
      p3_bit_slice_6574 <= p3_data_enable ? p2_bit_slice_6574 : p3_bit_slice_6574;
      p3_bit_slice_6575 <= p3_data_enable ? p2_bit_slice_6575 : p3_bit_slice_6575;
      p4_b <= p4_data_enable ? p3_b : p4_b;
      p4_uge_6652 <= p4_data_enable ? p3_uge_6652 : p4_uge_6652;
      p4_bivisor__1 <= p4_data_enable ? p3_bivisor__1 : p4_bivisor__1;
      p4_uge_6732 <= p4_data_enable ? p3_uge_6732 : p4_uge_6732;
      p4_uge_6810 <= p4_data_enable ? p3_uge_6810 : p4_uge_6810;
      p4_uge_6888 <= p4_data_enable ? uge_6888 : p4_uge_6888;
      p4_r__8 <= p4_data_enable ? r__8 : p4_r__8;
      p4_bit_slice_6548 <= p4_data_enable ? p3_bit_slice_6548 : p4_bit_slice_6548;
      p4_bit_slice_6549 <= p4_data_enable ? p3_bit_slice_6549 : p4_bit_slice_6549;
      p4_bit_slice_6550 <= p4_data_enable ? p3_bit_slice_6550 : p4_bit_slice_6550;
      p4_bit_slice_6551 <= p4_data_enable ? p3_bit_slice_6551 : p4_bit_slice_6551;
      p4_bit_slice_6552 <= p4_data_enable ? p3_bit_slice_6552 : p4_bit_slice_6552;
      p4_bit_slice_6553 <= p4_data_enable ? p3_bit_slice_6553 : p4_bit_slice_6553;
      p4_bit_slice_6554 <= p4_data_enable ? p3_bit_slice_6554 : p4_bit_slice_6554;
      p4_bit_slice_6555 <= p4_data_enable ? p3_bit_slice_6555 : p4_bit_slice_6555;
      p4_bit_slice_6556 <= p4_data_enable ? p3_bit_slice_6556 : p4_bit_slice_6556;
      p4_bit_slice_6557 <= p4_data_enable ? p3_bit_slice_6557 : p4_bit_slice_6557;
      p4_bit_slice_6558 <= p4_data_enable ? p3_bit_slice_6558 : p4_bit_slice_6558;
      p4_bit_slice_6559 <= p4_data_enable ? p3_bit_slice_6559 : p4_bit_slice_6559;
      p4_bit_slice_6560 <= p4_data_enable ? p3_bit_slice_6560 : p4_bit_slice_6560;
      p4_bit_slice_6561 <= p4_data_enable ? p3_bit_slice_6561 : p4_bit_slice_6561;
      p4_bit_slice_6562 <= p4_data_enable ? p3_bit_slice_6562 : p4_bit_slice_6562;
      p4_bit_slice_6563 <= p4_data_enable ? p3_bit_slice_6563 : p4_bit_slice_6563;
      p4_bit_slice_6564 <= p4_data_enable ? p3_bit_slice_6564 : p4_bit_slice_6564;
      p4_bit_slice_6565 <= p4_data_enable ? p3_bit_slice_6565 : p4_bit_slice_6565;
      p4_bit_slice_6566 <= p4_data_enable ? p3_bit_slice_6566 : p4_bit_slice_6566;
      p4_bit_slice_6567 <= p4_data_enable ? p3_bit_slice_6567 : p4_bit_slice_6567;
      p4_bit_slice_6568 <= p4_data_enable ? p3_bit_slice_6568 : p4_bit_slice_6568;
      p4_bit_slice_6569 <= p4_data_enable ? p3_bit_slice_6569 : p4_bit_slice_6569;
      p4_bit_slice_6570 <= p4_data_enable ? p3_bit_slice_6570 : p4_bit_slice_6570;
      p4_bit_slice_6571 <= p4_data_enable ? p3_bit_slice_6571 : p4_bit_slice_6571;
      p4_bit_slice_6572 <= p4_data_enable ? p3_bit_slice_6572 : p4_bit_slice_6572;
      p4_bit_slice_6573 <= p4_data_enable ? p3_bit_slice_6573 : p4_bit_slice_6573;
      p4_bit_slice_6574 <= p4_data_enable ? p3_bit_slice_6574 : p4_bit_slice_6574;
      p4_bit_slice_6575 <= p4_data_enable ? p3_bit_slice_6575 : p4_bit_slice_6575;
      p5_b <= p5_data_enable ? p4_b : p5_b;
      p5_uge_6652 <= p5_data_enable ? p4_uge_6652 : p5_uge_6652;
      p5_bivisor__1 <= p5_data_enable ? p4_bivisor__1 : p5_bivisor__1;
      p5_uge_6732 <= p5_data_enable ? p4_uge_6732 : p5_uge_6732;
      p5_uge_6810 <= p5_data_enable ? p4_uge_6810 : p5_uge_6810;
      p5_uge_6888 <= p5_data_enable ? p4_uge_6888 : p5_uge_6888;
      p5_uge_6966 <= p5_data_enable ? uge_6966 : p5_uge_6966;
      p5_r__10 <= p5_data_enable ? r__10 : p5_r__10;
      p5_bit_slice_6549 <= p5_data_enable ? p4_bit_slice_6549 : p5_bit_slice_6549;
      p5_bit_slice_6550 <= p5_data_enable ? p4_bit_slice_6550 : p5_bit_slice_6550;
      p5_bit_slice_6551 <= p5_data_enable ? p4_bit_slice_6551 : p5_bit_slice_6551;
      p5_bit_slice_6552 <= p5_data_enable ? p4_bit_slice_6552 : p5_bit_slice_6552;
      p5_bit_slice_6553 <= p5_data_enable ? p4_bit_slice_6553 : p5_bit_slice_6553;
      p5_bit_slice_6554 <= p5_data_enable ? p4_bit_slice_6554 : p5_bit_slice_6554;
      p5_bit_slice_6555 <= p5_data_enable ? p4_bit_slice_6555 : p5_bit_slice_6555;
      p5_bit_slice_6556 <= p5_data_enable ? p4_bit_slice_6556 : p5_bit_slice_6556;
      p5_bit_slice_6557 <= p5_data_enable ? p4_bit_slice_6557 : p5_bit_slice_6557;
      p5_bit_slice_6558 <= p5_data_enable ? p4_bit_slice_6558 : p5_bit_slice_6558;
      p5_bit_slice_6559 <= p5_data_enable ? p4_bit_slice_6559 : p5_bit_slice_6559;
      p5_bit_slice_6560 <= p5_data_enable ? p4_bit_slice_6560 : p5_bit_slice_6560;
      p5_bit_slice_6561 <= p5_data_enable ? p4_bit_slice_6561 : p5_bit_slice_6561;
      p5_bit_slice_6562 <= p5_data_enable ? p4_bit_slice_6562 : p5_bit_slice_6562;
      p5_bit_slice_6563 <= p5_data_enable ? p4_bit_slice_6563 : p5_bit_slice_6563;
      p5_bit_slice_6564 <= p5_data_enable ? p4_bit_slice_6564 : p5_bit_slice_6564;
      p5_bit_slice_6565 <= p5_data_enable ? p4_bit_slice_6565 : p5_bit_slice_6565;
      p5_bit_slice_6566 <= p5_data_enable ? p4_bit_slice_6566 : p5_bit_slice_6566;
      p5_bit_slice_6567 <= p5_data_enable ? p4_bit_slice_6567 : p5_bit_slice_6567;
      p5_bit_slice_6568 <= p5_data_enable ? p4_bit_slice_6568 : p5_bit_slice_6568;
      p5_bit_slice_6569 <= p5_data_enable ? p4_bit_slice_6569 : p5_bit_slice_6569;
      p5_bit_slice_6570 <= p5_data_enable ? p4_bit_slice_6570 : p5_bit_slice_6570;
      p5_bit_slice_6571 <= p5_data_enable ? p4_bit_slice_6571 : p5_bit_slice_6571;
      p5_bit_slice_6572 <= p5_data_enable ? p4_bit_slice_6572 : p5_bit_slice_6572;
      p5_bit_slice_6573 <= p5_data_enable ? p4_bit_slice_6573 : p5_bit_slice_6573;
      p5_bit_slice_6574 <= p5_data_enable ? p4_bit_slice_6574 : p5_bit_slice_6574;
      p5_bit_slice_6575 <= p5_data_enable ? p4_bit_slice_6575 : p5_bit_slice_6575;
      p6_b <= p6_data_enable ? p5_b : p6_b;
      p6_uge_6652 <= p6_data_enable ? p5_uge_6652 : p6_uge_6652;
      p6_bivisor__1 <= p6_data_enable ? p5_bivisor__1 : p6_bivisor__1;
      p6_uge_6732 <= p6_data_enable ? p5_uge_6732 : p6_uge_6732;
      p6_uge_6810 <= p6_data_enable ? p5_uge_6810 : p6_uge_6810;
      p6_uge_6888 <= p6_data_enable ? p5_uge_6888 : p6_uge_6888;
      p6_uge_6966 <= p6_data_enable ? p5_uge_6966 : p6_uge_6966;
      p6_uge_7044 <= p6_data_enable ? uge_7044 : p6_uge_7044;
      p6_r__12 <= p6_data_enable ? r__12 : p6_r__12;
      p6_bit_slice_6550 <= p6_data_enable ? p5_bit_slice_6550 : p6_bit_slice_6550;
      p6_bit_slice_6551 <= p6_data_enable ? p5_bit_slice_6551 : p6_bit_slice_6551;
      p6_bit_slice_6552 <= p6_data_enable ? p5_bit_slice_6552 : p6_bit_slice_6552;
      p6_bit_slice_6553 <= p6_data_enable ? p5_bit_slice_6553 : p6_bit_slice_6553;
      p6_bit_slice_6554 <= p6_data_enable ? p5_bit_slice_6554 : p6_bit_slice_6554;
      p6_bit_slice_6555 <= p6_data_enable ? p5_bit_slice_6555 : p6_bit_slice_6555;
      p6_bit_slice_6556 <= p6_data_enable ? p5_bit_slice_6556 : p6_bit_slice_6556;
      p6_bit_slice_6557 <= p6_data_enable ? p5_bit_slice_6557 : p6_bit_slice_6557;
      p6_bit_slice_6558 <= p6_data_enable ? p5_bit_slice_6558 : p6_bit_slice_6558;
      p6_bit_slice_6559 <= p6_data_enable ? p5_bit_slice_6559 : p6_bit_slice_6559;
      p6_bit_slice_6560 <= p6_data_enable ? p5_bit_slice_6560 : p6_bit_slice_6560;
      p6_bit_slice_6561 <= p6_data_enable ? p5_bit_slice_6561 : p6_bit_slice_6561;
      p6_bit_slice_6562 <= p6_data_enable ? p5_bit_slice_6562 : p6_bit_slice_6562;
      p6_bit_slice_6563 <= p6_data_enable ? p5_bit_slice_6563 : p6_bit_slice_6563;
      p6_bit_slice_6564 <= p6_data_enable ? p5_bit_slice_6564 : p6_bit_slice_6564;
      p6_bit_slice_6565 <= p6_data_enable ? p5_bit_slice_6565 : p6_bit_slice_6565;
      p6_bit_slice_6566 <= p6_data_enable ? p5_bit_slice_6566 : p6_bit_slice_6566;
      p6_bit_slice_6567 <= p6_data_enable ? p5_bit_slice_6567 : p6_bit_slice_6567;
      p6_bit_slice_6568 <= p6_data_enable ? p5_bit_slice_6568 : p6_bit_slice_6568;
      p6_bit_slice_6569 <= p6_data_enable ? p5_bit_slice_6569 : p6_bit_slice_6569;
      p6_bit_slice_6570 <= p6_data_enable ? p5_bit_slice_6570 : p6_bit_slice_6570;
      p6_bit_slice_6571 <= p6_data_enable ? p5_bit_slice_6571 : p6_bit_slice_6571;
      p6_bit_slice_6572 <= p6_data_enable ? p5_bit_slice_6572 : p6_bit_slice_6572;
      p6_bit_slice_6573 <= p6_data_enable ? p5_bit_slice_6573 : p6_bit_slice_6573;
      p6_bit_slice_6574 <= p6_data_enable ? p5_bit_slice_6574 : p6_bit_slice_6574;
      p6_bit_slice_6575 <= p6_data_enable ? p5_bit_slice_6575 : p6_bit_slice_6575;
      p7_b <= p7_data_enable ? p6_b : p7_b;
      p7_uge_6652 <= p7_data_enable ? p6_uge_6652 : p7_uge_6652;
      p7_bivisor__1 <= p7_data_enable ? p6_bivisor__1 : p7_bivisor__1;
      p7_uge_6732 <= p7_data_enable ? p6_uge_6732 : p7_uge_6732;
      p7_uge_6810 <= p7_data_enable ? p6_uge_6810 : p7_uge_6810;
      p7_uge_6888 <= p7_data_enable ? p6_uge_6888 : p7_uge_6888;
      p7_uge_6966 <= p7_data_enable ? p6_uge_6966 : p7_uge_6966;
      p7_uge_7044 <= p7_data_enable ? p6_uge_7044 : p7_uge_7044;
      p7_uge_7122 <= p7_data_enable ? uge_7122 : p7_uge_7122;
      p7_r__14 <= p7_data_enable ? r__14 : p7_r__14;
      p7_bit_slice_6551 <= p7_data_enable ? p6_bit_slice_6551 : p7_bit_slice_6551;
      p7_bit_slice_6552 <= p7_data_enable ? p6_bit_slice_6552 : p7_bit_slice_6552;
      p7_bit_slice_6553 <= p7_data_enable ? p6_bit_slice_6553 : p7_bit_slice_6553;
      p7_bit_slice_6554 <= p7_data_enable ? p6_bit_slice_6554 : p7_bit_slice_6554;
      p7_bit_slice_6555 <= p7_data_enable ? p6_bit_slice_6555 : p7_bit_slice_6555;
      p7_bit_slice_6556 <= p7_data_enable ? p6_bit_slice_6556 : p7_bit_slice_6556;
      p7_bit_slice_6557 <= p7_data_enable ? p6_bit_slice_6557 : p7_bit_slice_6557;
      p7_bit_slice_6558 <= p7_data_enable ? p6_bit_slice_6558 : p7_bit_slice_6558;
      p7_bit_slice_6559 <= p7_data_enable ? p6_bit_slice_6559 : p7_bit_slice_6559;
      p7_bit_slice_6560 <= p7_data_enable ? p6_bit_slice_6560 : p7_bit_slice_6560;
      p7_bit_slice_6561 <= p7_data_enable ? p6_bit_slice_6561 : p7_bit_slice_6561;
      p7_bit_slice_6562 <= p7_data_enable ? p6_bit_slice_6562 : p7_bit_slice_6562;
      p7_bit_slice_6563 <= p7_data_enable ? p6_bit_slice_6563 : p7_bit_slice_6563;
      p7_bit_slice_6564 <= p7_data_enable ? p6_bit_slice_6564 : p7_bit_slice_6564;
      p7_bit_slice_6565 <= p7_data_enable ? p6_bit_slice_6565 : p7_bit_slice_6565;
      p7_bit_slice_6566 <= p7_data_enable ? p6_bit_slice_6566 : p7_bit_slice_6566;
      p7_bit_slice_6567 <= p7_data_enable ? p6_bit_slice_6567 : p7_bit_slice_6567;
      p7_bit_slice_6568 <= p7_data_enable ? p6_bit_slice_6568 : p7_bit_slice_6568;
      p7_bit_slice_6569 <= p7_data_enable ? p6_bit_slice_6569 : p7_bit_slice_6569;
      p7_bit_slice_6570 <= p7_data_enable ? p6_bit_slice_6570 : p7_bit_slice_6570;
      p7_bit_slice_6571 <= p7_data_enable ? p6_bit_slice_6571 : p7_bit_slice_6571;
      p7_bit_slice_6572 <= p7_data_enable ? p6_bit_slice_6572 : p7_bit_slice_6572;
      p7_bit_slice_6573 <= p7_data_enable ? p6_bit_slice_6573 : p7_bit_slice_6573;
      p7_bit_slice_6574 <= p7_data_enable ? p6_bit_slice_6574 : p7_bit_slice_6574;
      p7_bit_slice_6575 <= p7_data_enable ? p6_bit_slice_6575 : p7_bit_slice_6575;
      p8_b <= p8_data_enable ? p7_b : p8_b;
      p8_uge_6652 <= p8_data_enable ? p7_uge_6652 : p8_uge_6652;
      p8_bivisor__1 <= p8_data_enable ? p7_bivisor__1 : p8_bivisor__1;
      p8_uge_6732 <= p8_data_enable ? p7_uge_6732 : p8_uge_6732;
      p8_uge_6810 <= p8_data_enable ? p7_uge_6810 : p8_uge_6810;
      p8_uge_6888 <= p8_data_enable ? p7_uge_6888 : p8_uge_6888;
      p8_uge_6966 <= p8_data_enable ? p7_uge_6966 : p8_uge_6966;
      p8_uge_7044 <= p8_data_enable ? p7_uge_7044 : p8_uge_7044;
      p8_uge_7122 <= p8_data_enable ? p7_uge_7122 : p8_uge_7122;
      p8_uge_7200 <= p8_data_enable ? uge_7200 : p8_uge_7200;
      p8_r__16 <= p8_data_enable ? r__16 : p8_r__16;
      p8_bit_slice_6552 <= p8_data_enable ? p7_bit_slice_6552 : p8_bit_slice_6552;
      p8_bit_slice_6553 <= p8_data_enable ? p7_bit_slice_6553 : p8_bit_slice_6553;
      p8_bit_slice_6554 <= p8_data_enable ? p7_bit_slice_6554 : p8_bit_slice_6554;
      p8_bit_slice_6555 <= p8_data_enable ? p7_bit_slice_6555 : p8_bit_slice_6555;
      p8_bit_slice_6556 <= p8_data_enable ? p7_bit_slice_6556 : p8_bit_slice_6556;
      p8_bit_slice_6557 <= p8_data_enable ? p7_bit_slice_6557 : p8_bit_slice_6557;
      p8_bit_slice_6558 <= p8_data_enable ? p7_bit_slice_6558 : p8_bit_slice_6558;
      p8_bit_slice_6559 <= p8_data_enable ? p7_bit_slice_6559 : p8_bit_slice_6559;
      p8_bit_slice_6560 <= p8_data_enable ? p7_bit_slice_6560 : p8_bit_slice_6560;
      p8_bit_slice_6561 <= p8_data_enable ? p7_bit_slice_6561 : p8_bit_slice_6561;
      p8_bit_slice_6562 <= p8_data_enable ? p7_bit_slice_6562 : p8_bit_slice_6562;
      p8_bit_slice_6563 <= p8_data_enable ? p7_bit_slice_6563 : p8_bit_slice_6563;
      p8_bit_slice_6564 <= p8_data_enable ? p7_bit_slice_6564 : p8_bit_slice_6564;
      p8_bit_slice_6565 <= p8_data_enable ? p7_bit_slice_6565 : p8_bit_slice_6565;
      p8_bit_slice_6566 <= p8_data_enable ? p7_bit_slice_6566 : p8_bit_slice_6566;
      p8_bit_slice_6567 <= p8_data_enable ? p7_bit_slice_6567 : p8_bit_slice_6567;
      p8_bit_slice_6568 <= p8_data_enable ? p7_bit_slice_6568 : p8_bit_slice_6568;
      p8_bit_slice_6569 <= p8_data_enable ? p7_bit_slice_6569 : p8_bit_slice_6569;
      p8_bit_slice_6570 <= p8_data_enable ? p7_bit_slice_6570 : p8_bit_slice_6570;
      p8_bit_slice_6571 <= p8_data_enable ? p7_bit_slice_6571 : p8_bit_slice_6571;
      p8_bit_slice_6572 <= p8_data_enable ? p7_bit_slice_6572 : p8_bit_slice_6572;
      p8_bit_slice_6573 <= p8_data_enable ? p7_bit_slice_6573 : p8_bit_slice_6573;
      p8_bit_slice_6574 <= p8_data_enable ? p7_bit_slice_6574 : p8_bit_slice_6574;
      p8_bit_slice_6575 <= p8_data_enable ? p7_bit_slice_6575 : p8_bit_slice_6575;
      p9_b <= p9_data_enable ? p8_b : p9_b;
      p9_uge_6652 <= p9_data_enable ? p8_uge_6652 : p9_uge_6652;
      p9_bivisor__1 <= p9_data_enable ? p8_bivisor__1 : p9_bivisor__1;
      p9_uge_6732 <= p9_data_enable ? p8_uge_6732 : p9_uge_6732;
      p9_uge_6810 <= p9_data_enable ? p8_uge_6810 : p9_uge_6810;
      p9_uge_6888 <= p9_data_enable ? p8_uge_6888 : p9_uge_6888;
      p9_uge_6966 <= p9_data_enable ? p8_uge_6966 : p9_uge_6966;
      p9_uge_7044 <= p9_data_enable ? p8_uge_7044 : p9_uge_7044;
      p9_uge_7122 <= p9_data_enable ? p8_uge_7122 : p9_uge_7122;
      p9_uge_7200 <= p9_data_enable ? p8_uge_7200 : p9_uge_7200;
      p9_uge_7278 <= p9_data_enable ? uge_7278 : p9_uge_7278;
      p9_r__18 <= p9_data_enable ? r__18 : p9_r__18;
      p9_bit_slice_6553 <= p9_data_enable ? p8_bit_slice_6553 : p9_bit_slice_6553;
      p9_bit_slice_6554 <= p9_data_enable ? p8_bit_slice_6554 : p9_bit_slice_6554;
      p9_bit_slice_6555 <= p9_data_enable ? p8_bit_slice_6555 : p9_bit_slice_6555;
      p9_bit_slice_6556 <= p9_data_enable ? p8_bit_slice_6556 : p9_bit_slice_6556;
      p9_bit_slice_6557 <= p9_data_enable ? p8_bit_slice_6557 : p9_bit_slice_6557;
      p9_bit_slice_6558 <= p9_data_enable ? p8_bit_slice_6558 : p9_bit_slice_6558;
      p9_bit_slice_6559 <= p9_data_enable ? p8_bit_slice_6559 : p9_bit_slice_6559;
      p9_bit_slice_6560 <= p9_data_enable ? p8_bit_slice_6560 : p9_bit_slice_6560;
      p9_bit_slice_6561 <= p9_data_enable ? p8_bit_slice_6561 : p9_bit_slice_6561;
      p9_bit_slice_6562 <= p9_data_enable ? p8_bit_slice_6562 : p9_bit_slice_6562;
      p9_bit_slice_6563 <= p9_data_enable ? p8_bit_slice_6563 : p9_bit_slice_6563;
      p9_bit_slice_6564 <= p9_data_enable ? p8_bit_slice_6564 : p9_bit_slice_6564;
      p9_bit_slice_6565 <= p9_data_enable ? p8_bit_slice_6565 : p9_bit_slice_6565;
      p9_bit_slice_6566 <= p9_data_enable ? p8_bit_slice_6566 : p9_bit_slice_6566;
      p9_bit_slice_6567 <= p9_data_enable ? p8_bit_slice_6567 : p9_bit_slice_6567;
      p9_bit_slice_6568 <= p9_data_enable ? p8_bit_slice_6568 : p9_bit_slice_6568;
      p9_bit_slice_6569 <= p9_data_enable ? p8_bit_slice_6569 : p9_bit_slice_6569;
      p9_bit_slice_6570 <= p9_data_enable ? p8_bit_slice_6570 : p9_bit_slice_6570;
      p9_bit_slice_6571 <= p9_data_enable ? p8_bit_slice_6571 : p9_bit_slice_6571;
      p9_bit_slice_6572 <= p9_data_enable ? p8_bit_slice_6572 : p9_bit_slice_6572;
      p9_bit_slice_6573 <= p9_data_enable ? p8_bit_slice_6573 : p9_bit_slice_6573;
      p9_bit_slice_6574 <= p9_data_enable ? p8_bit_slice_6574 : p9_bit_slice_6574;
      p9_bit_slice_6575 <= p9_data_enable ? p8_bit_slice_6575 : p9_bit_slice_6575;
      p10_b <= p10_data_enable ? p9_b : p10_b;
      p10_uge_6652 <= p10_data_enable ? p9_uge_6652 : p10_uge_6652;
      p10_bivisor__1 <= p10_data_enable ? p9_bivisor__1 : p10_bivisor__1;
      p10_uge_6732 <= p10_data_enable ? p9_uge_6732 : p10_uge_6732;
      p10_uge_6810 <= p10_data_enable ? p9_uge_6810 : p10_uge_6810;
      p10_uge_6888 <= p10_data_enable ? p9_uge_6888 : p10_uge_6888;
      p10_uge_6966 <= p10_data_enable ? p9_uge_6966 : p10_uge_6966;
      p10_uge_7044 <= p10_data_enable ? p9_uge_7044 : p10_uge_7044;
      p10_uge_7122 <= p10_data_enable ? p9_uge_7122 : p10_uge_7122;
      p10_uge_7200 <= p10_data_enable ? p9_uge_7200 : p10_uge_7200;
      p10_uge_7278 <= p10_data_enable ? p9_uge_7278 : p10_uge_7278;
      p10_uge_7356 <= p10_data_enable ? uge_7356 : p10_uge_7356;
      p10_r__20 <= p10_data_enable ? r__20 : p10_r__20;
      p10_bit_slice_6554 <= p10_data_enable ? p9_bit_slice_6554 : p10_bit_slice_6554;
      p10_bit_slice_6555 <= p10_data_enable ? p9_bit_slice_6555 : p10_bit_slice_6555;
      p10_bit_slice_6556 <= p10_data_enable ? p9_bit_slice_6556 : p10_bit_slice_6556;
      p10_bit_slice_6557 <= p10_data_enable ? p9_bit_slice_6557 : p10_bit_slice_6557;
      p10_bit_slice_6558 <= p10_data_enable ? p9_bit_slice_6558 : p10_bit_slice_6558;
      p10_bit_slice_6559 <= p10_data_enable ? p9_bit_slice_6559 : p10_bit_slice_6559;
      p10_bit_slice_6560 <= p10_data_enable ? p9_bit_slice_6560 : p10_bit_slice_6560;
      p10_bit_slice_6561 <= p10_data_enable ? p9_bit_slice_6561 : p10_bit_slice_6561;
      p10_bit_slice_6562 <= p10_data_enable ? p9_bit_slice_6562 : p10_bit_slice_6562;
      p10_bit_slice_6563 <= p10_data_enable ? p9_bit_slice_6563 : p10_bit_slice_6563;
      p10_bit_slice_6564 <= p10_data_enable ? p9_bit_slice_6564 : p10_bit_slice_6564;
      p10_bit_slice_6565 <= p10_data_enable ? p9_bit_slice_6565 : p10_bit_slice_6565;
      p10_bit_slice_6566 <= p10_data_enable ? p9_bit_slice_6566 : p10_bit_slice_6566;
      p10_bit_slice_6567 <= p10_data_enable ? p9_bit_slice_6567 : p10_bit_slice_6567;
      p10_bit_slice_6568 <= p10_data_enable ? p9_bit_slice_6568 : p10_bit_slice_6568;
      p10_bit_slice_6569 <= p10_data_enable ? p9_bit_slice_6569 : p10_bit_slice_6569;
      p10_bit_slice_6570 <= p10_data_enable ? p9_bit_slice_6570 : p10_bit_slice_6570;
      p10_bit_slice_6571 <= p10_data_enable ? p9_bit_slice_6571 : p10_bit_slice_6571;
      p10_bit_slice_6572 <= p10_data_enable ? p9_bit_slice_6572 : p10_bit_slice_6572;
      p10_bit_slice_6573 <= p10_data_enable ? p9_bit_slice_6573 : p10_bit_slice_6573;
      p10_bit_slice_6574 <= p10_data_enable ? p9_bit_slice_6574 : p10_bit_slice_6574;
      p10_bit_slice_6575 <= p10_data_enable ? p9_bit_slice_6575 : p10_bit_slice_6575;
      p11_b <= p11_data_enable ? p10_b : p11_b;
      p11_uge_6652 <= p11_data_enable ? p10_uge_6652 : p11_uge_6652;
      p11_bivisor__1 <= p11_data_enable ? p10_bivisor__1 : p11_bivisor__1;
      p11_uge_6732 <= p11_data_enable ? p10_uge_6732 : p11_uge_6732;
      p11_uge_6810 <= p11_data_enable ? p10_uge_6810 : p11_uge_6810;
      p11_uge_6888 <= p11_data_enable ? p10_uge_6888 : p11_uge_6888;
      p11_uge_6966 <= p11_data_enable ? p10_uge_6966 : p11_uge_6966;
      p11_uge_7044 <= p11_data_enable ? p10_uge_7044 : p11_uge_7044;
      p11_uge_7122 <= p11_data_enable ? p10_uge_7122 : p11_uge_7122;
      p11_uge_7200 <= p11_data_enable ? p10_uge_7200 : p11_uge_7200;
      p11_uge_7278 <= p11_data_enable ? p10_uge_7278 : p11_uge_7278;
      p11_uge_7356 <= p11_data_enable ? p10_uge_7356 : p11_uge_7356;
      p11_uge_7434 <= p11_data_enable ? uge_7434 : p11_uge_7434;
      p11_r__22 <= p11_data_enable ? r__22 : p11_r__22;
      p11_bit_slice_6555 <= p11_data_enable ? p10_bit_slice_6555 : p11_bit_slice_6555;
      p11_bit_slice_6556 <= p11_data_enable ? p10_bit_slice_6556 : p11_bit_slice_6556;
      p11_bit_slice_6557 <= p11_data_enable ? p10_bit_slice_6557 : p11_bit_slice_6557;
      p11_bit_slice_6558 <= p11_data_enable ? p10_bit_slice_6558 : p11_bit_slice_6558;
      p11_bit_slice_6559 <= p11_data_enable ? p10_bit_slice_6559 : p11_bit_slice_6559;
      p11_bit_slice_6560 <= p11_data_enable ? p10_bit_slice_6560 : p11_bit_slice_6560;
      p11_bit_slice_6561 <= p11_data_enable ? p10_bit_slice_6561 : p11_bit_slice_6561;
      p11_bit_slice_6562 <= p11_data_enable ? p10_bit_slice_6562 : p11_bit_slice_6562;
      p11_bit_slice_6563 <= p11_data_enable ? p10_bit_slice_6563 : p11_bit_slice_6563;
      p11_bit_slice_6564 <= p11_data_enable ? p10_bit_slice_6564 : p11_bit_slice_6564;
      p11_bit_slice_6565 <= p11_data_enable ? p10_bit_slice_6565 : p11_bit_slice_6565;
      p11_bit_slice_6566 <= p11_data_enable ? p10_bit_slice_6566 : p11_bit_slice_6566;
      p11_bit_slice_6567 <= p11_data_enable ? p10_bit_slice_6567 : p11_bit_slice_6567;
      p11_bit_slice_6568 <= p11_data_enable ? p10_bit_slice_6568 : p11_bit_slice_6568;
      p11_bit_slice_6569 <= p11_data_enable ? p10_bit_slice_6569 : p11_bit_slice_6569;
      p11_bit_slice_6570 <= p11_data_enable ? p10_bit_slice_6570 : p11_bit_slice_6570;
      p11_bit_slice_6571 <= p11_data_enable ? p10_bit_slice_6571 : p11_bit_slice_6571;
      p11_bit_slice_6572 <= p11_data_enable ? p10_bit_slice_6572 : p11_bit_slice_6572;
      p11_bit_slice_6573 <= p11_data_enable ? p10_bit_slice_6573 : p11_bit_slice_6573;
      p11_bit_slice_6574 <= p11_data_enable ? p10_bit_slice_6574 : p11_bit_slice_6574;
      p11_bit_slice_6575 <= p11_data_enable ? p10_bit_slice_6575 : p11_bit_slice_6575;
      p12_b <= p12_data_enable ? p11_b : p12_b;
      p12_uge_6652 <= p12_data_enable ? p11_uge_6652 : p12_uge_6652;
      p12_bivisor__1 <= p12_data_enable ? p11_bivisor__1 : p12_bivisor__1;
      p12_uge_6732 <= p12_data_enable ? p11_uge_6732 : p12_uge_6732;
      p12_uge_6810 <= p12_data_enable ? p11_uge_6810 : p12_uge_6810;
      p12_uge_6888 <= p12_data_enable ? p11_uge_6888 : p12_uge_6888;
      p12_uge_6966 <= p12_data_enable ? p11_uge_6966 : p12_uge_6966;
      p12_uge_7044 <= p12_data_enable ? p11_uge_7044 : p12_uge_7044;
      p12_uge_7122 <= p12_data_enable ? p11_uge_7122 : p12_uge_7122;
      p12_uge_7200 <= p12_data_enable ? p11_uge_7200 : p12_uge_7200;
      p12_uge_7278 <= p12_data_enable ? p11_uge_7278 : p12_uge_7278;
      p12_uge_7356 <= p12_data_enable ? p11_uge_7356 : p12_uge_7356;
      p12_uge_7434 <= p12_data_enable ? p11_uge_7434 : p12_uge_7434;
      p12_uge_7512 <= p12_data_enable ? uge_7512 : p12_uge_7512;
      p12_r__24 <= p12_data_enable ? r__24 : p12_r__24;
      p12_bit_slice_6556 <= p12_data_enable ? p11_bit_slice_6556 : p12_bit_slice_6556;
      p12_bit_slice_6557 <= p12_data_enable ? p11_bit_slice_6557 : p12_bit_slice_6557;
      p12_bit_slice_6558 <= p12_data_enable ? p11_bit_slice_6558 : p12_bit_slice_6558;
      p12_bit_slice_6559 <= p12_data_enable ? p11_bit_slice_6559 : p12_bit_slice_6559;
      p12_bit_slice_6560 <= p12_data_enable ? p11_bit_slice_6560 : p12_bit_slice_6560;
      p12_bit_slice_6561 <= p12_data_enable ? p11_bit_slice_6561 : p12_bit_slice_6561;
      p12_bit_slice_6562 <= p12_data_enable ? p11_bit_slice_6562 : p12_bit_slice_6562;
      p12_bit_slice_6563 <= p12_data_enable ? p11_bit_slice_6563 : p12_bit_slice_6563;
      p12_bit_slice_6564 <= p12_data_enable ? p11_bit_slice_6564 : p12_bit_slice_6564;
      p12_bit_slice_6565 <= p12_data_enable ? p11_bit_slice_6565 : p12_bit_slice_6565;
      p12_bit_slice_6566 <= p12_data_enable ? p11_bit_slice_6566 : p12_bit_slice_6566;
      p12_bit_slice_6567 <= p12_data_enable ? p11_bit_slice_6567 : p12_bit_slice_6567;
      p12_bit_slice_6568 <= p12_data_enable ? p11_bit_slice_6568 : p12_bit_slice_6568;
      p12_bit_slice_6569 <= p12_data_enable ? p11_bit_slice_6569 : p12_bit_slice_6569;
      p12_bit_slice_6570 <= p12_data_enable ? p11_bit_slice_6570 : p12_bit_slice_6570;
      p12_bit_slice_6571 <= p12_data_enable ? p11_bit_slice_6571 : p12_bit_slice_6571;
      p12_bit_slice_6572 <= p12_data_enable ? p11_bit_slice_6572 : p12_bit_slice_6572;
      p12_bit_slice_6573 <= p12_data_enable ? p11_bit_slice_6573 : p12_bit_slice_6573;
      p12_bit_slice_6574 <= p12_data_enable ? p11_bit_slice_6574 : p12_bit_slice_6574;
      p12_bit_slice_6575 <= p12_data_enable ? p11_bit_slice_6575 : p12_bit_slice_6575;
      p13_b <= p13_data_enable ? p12_b : p13_b;
      p13_uge_6652 <= p13_data_enable ? p12_uge_6652 : p13_uge_6652;
      p13_bivisor__1 <= p13_data_enable ? p12_bivisor__1 : p13_bivisor__1;
      p13_uge_6732 <= p13_data_enable ? p12_uge_6732 : p13_uge_6732;
      p13_uge_6810 <= p13_data_enable ? p12_uge_6810 : p13_uge_6810;
      p13_uge_6888 <= p13_data_enable ? p12_uge_6888 : p13_uge_6888;
      p13_uge_6966 <= p13_data_enable ? p12_uge_6966 : p13_uge_6966;
      p13_uge_7044 <= p13_data_enable ? p12_uge_7044 : p13_uge_7044;
      p13_uge_7122 <= p13_data_enable ? p12_uge_7122 : p13_uge_7122;
      p13_uge_7200 <= p13_data_enable ? p12_uge_7200 : p13_uge_7200;
      p13_uge_7278 <= p13_data_enable ? p12_uge_7278 : p13_uge_7278;
      p13_uge_7356 <= p13_data_enable ? p12_uge_7356 : p13_uge_7356;
      p13_uge_7434 <= p13_data_enable ? p12_uge_7434 : p13_uge_7434;
      p13_uge_7512 <= p13_data_enable ? p12_uge_7512 : p13_uge_7512;
      p13_uge_7590 <= p13_data_enable ? uge_7590 : p13_uge_7590;
      p13_r__26 <= p13_data_enable ? r__26 : p13_r__26;
      p13_bit_slice_6557 <= p13_data_enable ? p12_bit_slice_6557 : p13_bit_slice_6557;
      p13_bit_slice_6558 <= p13_data_enable ? p12_bit_slice_6558 : p13_bit_slice_6558;
      p13_bit_slice_6559 <= p13_data_enable ? p12_bit_slice_6559 : p13_bit_slice_6559;
      p13_bit_slice_6560 <= p13_data_enable ? p12_bit_slice_6560 : p13_bit_slice_6560;
      p13_bit_slice_6561 <= p13_data_enable ? p12_bit_slice_6561 : p13_bit_slice_6561;
      p13_bit_slice_6562 <= p13_data_enable ? p12_bit_slice_6562 : p13_bit_slice_6562;
      p13_bit_slice_6563 <= p13_data_enable ? p12_bit_slice_6563 : p13_bit_slice_6563;
      p13_bit_slice_6564 <= p13_data_enable ? p12_bit_slice_6564 : p13_bit_slice_6564;
      p13_bit_slice_6565 <= p13_data_enable ? p12_bit_slice_6565 : p13_bit_slice_6565;
      p13_bit_slice_6566 <= p13_data_enable ? p12_bit_slice_6566 : p13_bit_slice_6566;
      p13_bit_slice_6567 <= p13_data_enable ? p12_bit_slice_6567 : p13_bit_slice_6567;
      p13_bit_slice_6568 <= p13_data_enable ? p12_bit_slice_6568 : p13_bit_slice_6568;
      p13_bit_slice_6569 <= p13_data_enable ? p12_bit_slice_6569 : p13_bit_slice_6569;
      p13_bit_slice_6570 <= p13_data_enable ? p12_bit_slice_6570 : p13_bit_slice_6570;
      p13_bit_slice_6571 <= p13_data_enable ? p12_bit_slice_6571 : p13_bit_slice_6571;
      p13_bit_slice_6572 <= p13_data_enable ? p12_bit_slice_6572 : p13_bit_slice_6572;
      p13_bit_slice_6573 <= p13_data_enable ? p12_bit_slice_6573 : p13_bit_slice_6573;
      p13_bit_slice_6574 <= p13_data_enable ? p12_bit_slice_6574 : p13_bit_slice_6574;
      p13_bit_slice_6575 <= p13_data_enable ? p12_bit_slice_6575 : p13_bit_slice_6575;
      p14_b <= p14_data_enable ? p13_b : p14_b;
      p14_uge_6652 <= p14_data_enable ? p13_uge_6652 : p14_uge_6652;
      p14_bivisor__1 <= p14_data_enable ? p13_bivisor__1 : p14_bivisor__1;
      p14_uge_6732 <= p14_data_enable ? p13_uge_6732 : p14_uge_6732;
      p14_uge_6810 <= p14_data_enable ? p13_uge_6810 : p14_uge_6810;
      p14_uge_6888 <= p14_data_enable ? p13_uge_6888 : p14_uge_6888;
      p14_uge_6966 <= p14_data_enable ? p13_uge_6966 : p14_uge_6966;
      p14_uge_7044 <= p14_data_enable ? p13_uge_7044 : p14_uge_7044;
      p14_uge_7122 <= p14_data_enable ? p13_uge_7122 : p14_uge_7122;
      p14_uge_7200 <= p14_data_enable ? p13_uge_7200 : p14_uge_7200;
      p14_uge_7278 <= p14_data_enable ? p13_uge_7278 : p14_uge_7278;
      p14_uge_7356 <= p14_data_enable ? p13_uge_7356 : p14_uge_7356;
      p14_uge_7434 <= p14_data_enable ? p13_uge_7434 : p14_uge_7434;
      p14_uge_7512 <= p14_data_enable ? p13_uge_7512 : p14_uge_7512;
      p14_uge_7590 <= p14_data_enable ? p13_uge_7590 : p14_uge_7590;
      p14_uge_7668 <= p14_data_enable ? uge_7668 : p14_uge_7668;
      p14_r__28 <= p14_data_enable ? r__28 : p14_r__28;
      p14_bit_slice_6558 <= p14_data_enable ? p13_bit_slice_6558 : p14_bit_slice_6558;
      p14_bit_slice_6559 <= p14_data_enable ? p13_bit_slice_6559 : p14_bit_slice_6559;
      p14_bit_slice_6560 <= p14_data_enable ? p13_bit_slice_6560 : p14_bit_slice_6560;
      p14_bit_slice_6561 <= p14_data_enable ? p13_bit_slice_6561 : p14_bit_slice_6561;
      p14_bit_slice_6562 <= p14_data_enable ? p13_bit_slice_6562 : p14_bit_slice_6562;
      p14_bit_slice_6563 <= p14_data_enable ? p13_bit_slice_6563 : p14_bit_slice_6563;
      p14_bit_slice_6564 <= p14_data_enable ? p13_bit_slice_6564 : p14_bit_slice_6564;
      p14_bit_slice_6565 <= p14_data_enable ? p13_bit_slice_6565 : p14_bit_slice_6565;
      p14_bit_slice_6566 <= p14_data_enable ? p13_bit_slice_6566 : p14_bit_slice_6566;
      p14_bit_slice_6567 <= p14_data_enable ? p13_bit_slice_6567 : p14_bit_slice_6567;
      p14_bit_slice_6568 <= p14_data_enable ? p13_bit_slice_6568 : p14_bit_slice_6568;
      p14_bit_slice_6569 <= p14_data_enable ? p13_bit_slice_6569 : p14_bit_slice_6569;
      p14_bit_slice_6570 <= p14_data_enable ? p13_bit_slice_6570 : p14_bit_slice_6570;
      p14_bit_slice_6571 <= p14_data_enable ? p13_bit_slice_6571 : p14_bit_slice_6571;
      p14_bit_slice_6572 <= p14_data_enable ? p13_bit_slice_6572 : p14_bit_slice_6572;
      p14_bit_slice_6573 <= p14_data_enable ? p13_bit_slice_6573 : p14_bit_slice_6573;
      p14_bit_slice_6574 <= p14_data_enable ? p13_bit_slice_6574 : p14_bit_slice_6574;
      p14_bit_slice_6575 <= p14_data_enable ? p13_bit_slice_6575 : p14_bit_slice_6575;
      p15_b <= p15_data_enable ? p14_b : p15_b;
      p15_uge_6652 <= p15_data_enable ? p14_uge_6652 : p15_uge_6652;
      p15_bivisor__1 <= p15_data_enable ? p14_bivisor__1 : p15_bivisor__1;
      p15_uge_6732 <= p15_data_enable ? p14_uge_6732 : p15_uge_6732;
      p15_uge_6810 <= p15_data_enable ? p14_uge_6810 : p15_uge_6810;
      p15_uge_6888 <= p15_data_enable ? p14_uge_6888 : p15_uge_6888;
      p15_uge_6966 <= p15_data_enable ? p14_uge_6966 : p15_uge_6966;
      p15_uge_7044 <= p15_data_enable ? p14_uge_7044 : p15_uge_7044;
      p15_uge_7122 <= p15_data_enable ? p14_uge_7122 : p15_uge_7122;
      p15_uge_7200 <= p15_data_enable ? p14_uge_7200 : p15_uge_7200;
      p15_uge_7278 <= p15_data_enable ? p14_uge_7278 : p15_uge_7278;
      p15_uge_7356 <= p15_data_enable ? p14_uge_7356 : p15_uge_7356;
      p15_uge_7434 <= p15_data_enable ? p14_uge_7434 : p15_uge_7434;
      p15_uge_7512 <= p15_data_enable ? p14_uge_7512 : p15_uge_7512;
      p15_uge_7590 <= p15_data_enable ? p14_uge_7590 : p15_uge_7590;
      p15_uge_7668 <= p15_data_enable ? p14_uge_7668 : p15_uge_7668;
      p15_uge_7746 <= p15_data_enable ? uge_7746 : p15_uge_7746;
      p15_r__30 <= p15_data_enable ? r__30 : p15_r__30;
      p15_bit_slice_6559 <= p15_data_enable ? p14_bit_slice_6559 : p15_bit_slice_6559;
      p15_bit_slice_6560 <= p15_data_enable ? p14_bit_slice_6560 : p15_bit_slice_6560;
      p15_bit_slice_6561 <= p15_data_enable ? p14_bit_slice_6561 : p15_bit_slice_6561;
      p15_bit_slice_6562 <= p15_data_enable ? p14_bit_slice_6562 : p15_bit_slice_6562;
      p15_bit_slice_6563 <= p15_data_enable ? p14_bit_slice_6563 : p15_bit_slice_6563;
      p15_bit_slice_6564 <= p15_data_enable ? p14_bit_slice_6564 : p15_bit_slice_6564;
      p15_bit_slice_6565 <= p15_data_enable ? p14_bit_slice_6565 : p15_bit_slice_6565;
      p15_bit_slice_6566 <= p15_data_enable ? p14_bit_slice_6566 : p15_bit_slice_6566;
      p15_bit_slice_6567 <= p15_data_enable ? p14_bit_slice_6567 : p15_bit_slice_6567;
      p15_bit_slice_6568 <= p15_data_enable ? p14_bit_slice_6568 : p15_bit_slice_6568;
      p15_bit_slice_6569 <= p15_data_enable ? p14_bit_slice_6569 : p15_bit_slice_6569;
      p15_bit_slice_6570 <= p15_data_enable ? p14_bit_slice_6570 : p15_bit_slice_6570;
      p15_bit_slice_6571 <= p15_data_enable ? p14_bit_slice_6571 : p15_bit_slice_6571;
      p15_bit_slice_6572 <= p15_data_enable ? p14_bit_slice_6572 : p15_bit_slice_6572;
      p15_bit_slice_6573 <= p15_data_enable ? p14_bit_slice_6573 : p15_bit_slice_6573;
      p15_bit_slice_6574 <= p15_data_enable ? p14_bit_slice_6574 : p15_bit_slice_6574;
      p15_bit_slice_6575 <= p15_data_enable ? p14_bit_slice_6575 : p15_bit_slice_6575;
      p16_b <= p16_data_enable ? p15_b : p16_b;
      p16_uge_6652 <= p16_data_enable ? p15_uge_6652 : p16_uge_6652;
      p16_bivisor__1 <= p16_data_enable ? p15_bivisor__1 : p16_bivisor__1;
      p16_uge_6732 <= p16_data_enable ? p15_uge_6732 : p16_uge_6732;
      p16_uge_6810 <= p16_data_enable ? p15_uge_6810 : p16_uge_6810;
      p16_uge_6888 <= p16_data_enable ? p15_uge_6888 : p16_uge_6888;
      p16_uge_6966 <= p16_data_enable ? p15_uge_6966 : p16_uge_6966;
      p16_uge_7044 <= p16_data_enable ? p15_uge_7044 : p16_uge_7044;
      p16_uge_7122 <= p16_data_enable ? p15_uge_7122 : p16_uge_7122;
      p16_uge_7200 <= p16_data_enable ? p15_uge_7200 : p16_uge_7200;
      p16_uge_7278 <= p16_data_enable ? p15_uge_7278 : p16_uge_7278;
      p16_uge_7356 <= p16_data_enable ? p15_uge_7356 : p16_uge_7356;
      p16_uge_7434 <= p16_data_enable ? p15_uge_7434 : p16_uge_7434;
      p16_uge_7512 <= p16_data_enable ? p15_uge_7512 : p16_uge_7512;
      p16_uge_7590 <= p16_data_enable ? p15_uge_7590 : p16_uge_7590;
      p16_uge_7668 <= p16_data_enable ? p15_uge_7668 : p16_uge_7668;
      p16_uge_7746 <= p16_data_enable ? p15_uge_7746 : p16_uge_7746;
      p16_uge_7824 <= p16_data_enable ? uge_7824 : p16_uge_7824;
      p16_r__32 <= p16_data_enable ? r__32 : p16_r__32;
      p16_bit_slice_6560 <= p16_data_enable ? p15_bit_slice_6560 : p16_bit_slice_6560;
      p16_bit_slice_6561 <= p16_data_enable ? p15_bit_slice_6561 : p16_bit_slice_6561;
      p16_bit_slice_6562 <= p16_data_enable ? p15_bit_slice_6562 : p16_bit_slice_6562;
      p16_bit_slice_6563 <= p16_data_enable ? p15_bit_slice_6563 : p16_bit_slice_6563;
      p16_bit_slice_6564 <= p16_data_enable ? p15_bit_slice_6564 : p16_bit_slice_6564;
      p16_bit_slice_6565 <= p16_data_enable ? p15_bit_slice_6565 : p16_bit_slice_6565;
      p16_bit_slice_6566 <= p16_data_enable ? p15_bit_slice_6566 : p16_bit_slice_6566;
      p16_bit_slice_6567 <= p16_data_enable ? p15_bit_slice_6567 : p16_bit_slice_6567;
      p16_bit_slice_6568 <= p16_data_enable ? p15_bit_slice_6568 : p16_bit_slice_6568;
      p16_bit_slice_6569 <= p16_data_enable ? p15_bit_slice_6569 : p16_bit_slice_6569;
      p16_bit_slice_6570 <= p16_data_enable ? p15_bit_slice_6570 : p16_bit_slice_6570;
      p16_bit_slice_6571 <= p16_data_enable ? p15_bit_slice_6571 : p16_bit_slice_6571;
      p16_bit_slice_6572 <= p16_data_enable ? p15_bit_slice_6572 : p16_bit_slice_6572;
      p16_bit_slice_6573 <= p16_data_enable ? p15_bit_slice_6573 : p16_bit_slice_6573;
      p16_bit_slice_6574 <= p16_data_enable ? p15_bit_slice_6574 : p16_bit_slice_6574;
      p16_bit_slice_6575 <= p16_data_enable ? p15_bit_slice_6575 : p16_bit_slice_6575;
      p17_b <= p17_data_enable ? p16_b : p17_b;
      p17_uge_6652 <= p17_data_enable ? p16_uge_6652 : p17_uge_6652;
      p17_bivisor__1 <= p17_data_enable ? p16_bivisor__1 : p17_bivisor__1;
      p17_uge_6732 <= p17_data_enable ? p16_uge_6732 : p17_uge_6732;
      p17_uge_6810 <= p17_data_enable ? p16_uge_6810 : p17_uge_6810;
      p17_uge_6888 <= p17_data_enable ? p16_uge_6888 : p17_uge_6888;
      p17_uge_6966 <= p17_data_enable ? p16_uge_6966 : p17_uge_6966;
      p17_uge_7044 <= p17_data_enable ? p16_uge_7044 : p17_uge_7044;
      p17_uge_7122 <= p17_data_enable ? p16_uge_7122 : p17_uge_7122;
      p17_uge_7200 <= p17_data_enable ? p16_uge_7200 : p17_uge_7200;
      p17_uge_7278 <= p17_data_enable ? p16_uge_7278 : p17_uge_7278;
      p17_uge_7356 <= p17_data_enable ? p16_uge_7356 : p17_uge_7356;
      p17_uge_7434 <= p17_data_enable ? p16_uge_7434 : p17_uge_7434;
      p17_uge_7512 <= p17_data_enable ? p16_uge_7512 : p17_uge_7512;
      p17_uge_7590 <= p17_data_enable ? p16_uge_7590 : p17_uge_7590;
      p17_uge_7668 <= p17_data_enable ? p16_uge_7668 : p17_uge_7668;
      p17_uge_7746 <= p17_data_enable ? p16_uge_7746 : p17_uge_7746;
      p17_uge_7824 <= p17_data_enable ? p16_uge_7824 : p17_uge_7824;
      p17_uge_7902 <= p17_data_enable ? uge_7902 : p17_uge_7902;
      p17_r__34 <= p17_data_enable ? r__34 : p17_r__34;
      p17_bit_slice_6561 <= p17_data_enable ? p16_bit_slice_6561 : p17_bit_slice_6561;
      p17_bit_slice_6562 <= p17_data_enable ? p16_bit_slice_6562 : p17_bit_slice_6562;
      p17_bit_slice_6563 <= p17_data_enable ? p16_bit_slice_6563 : p17_bit_slice_6563;
      p17_bit_slice_6564 <= p17_data_enable ? p16_bit_slice_6564 : p17_bit_slice_6564;
      p17_bit_slice_6565 <= p17_data_enable ? p16_bit_slice_6565 : p17_bit_slice_6565;
      p17_bit_slice_6566 <= p17_data_enable ? p16_bit_slice_6566 : p17_bit_slice_6566;
      p17_bit_slice_6567 <= p17_data_enable ? p16_bit_slice_6567 : p17_bit_slice_6567;
      p17_bit_slice_6568 <= p17_data_enable ? p16_bit_slice_6568 : p17_bit_slice_6568;
      p17_bit_slice_6569 <= p17_data_enable ? p16_bit_slice_6569 : p17_bit_slice_6569;
      p17_bit_slice_6570 <= p17_data_enable ? p16_bit_slice_6570 : p17_bit_slice_6570;
      p17_bit_slice_6571 <= p17_data_enable ? p16_bit_slice_6571 : p17_bit_slice_6571;
      p17_bit_slice_6572 <= p17_data_enable ? p16_bit_slice_6572 : p17_bit_slice_6572;
      p17_bit_slice_6573 <= p17_data_enable ? p16_bit_slice_6573 : p17_bit_slice_6573;
      p17_bit_slice_6574 <= p17_data_enable ? p16_bit_slice_6574 : p17_bit_slice_6574;
      p17_bit_slice_6575 <= p17_data_enable ? p16_bit_slice_6575 : p17_bit_slice_6575;
      p18_b <= p18_data_enable ? p17_b : p18_b;
      p18_uge_6652 <= p18_data_enable ? p17_uge_6652 : p18_uge_6652;
      p18_bivisor__1 <= p18_data_enable ? p17_bivisor__1 : p18_bivisor__1;
      p18_uge_6732 <= p18_data_enable ? p17_uge_6732 : p18_uge_6732;
      p18_uge_6810 <= p18_data_enable ? p17_uge_6810 : p18_uge_6810;
      p18_uge_6888 <= p18_data_enable ? p17_uge_6888 : p18_uge_6888;
      p18_uge_6966 <= p18_data_enable ? p17_uge_6966 : p18_uge_6966;
      p18_uge_7044 <= p18_data_enable ? p17_uge_7044 : p18_uge_7044;
      p18_uge_7122 <= p18_data_enable ? p17_uge_7122 : p18_uge_7122;
      p18_uge_7200 <= p18_data_enable ? p17_uge_7200 : p18_uge_7200;
      p18_uge_7278 <= p18_data_enable ? p17_uge_7278 : p18_uge_7278;
      p18_uge_7356 <= p18_data_enable ? p17_uge_7356 : p18_uge_7356;
      p18_uge_7434 <= p18_data_enable ? p17_uge_7434 : p18_uge_7434;
      p18_uge_7512 <= p18_data_enable ? p17_uge_7512 : p18_uge_7512;
      p18_uge_7590 <= p18_data_enable ? p17_uge_7590 : p18_uge_7590;
      p18_uge_7668 <= p18_data_enable ? p17_uge_7668 : p18_uge_7668;
      p18_uge_7746 <= p18_data_enable ? p17_uge_7746 : p18_uge_7746;
      p18_uge_7824 <= p18_data_enable ? p17_uge_7824 : p18_uge_7824;
      p18_uge_7902 <= p18_data_enable ? p17_uge_7902 : p18_uge_7902;
      p18_uge_7980 <= p18_data_enable ? uge_7980 : p18_uge_7980;
      p18_r__36 <= p18_data_enable ? r__36 : p18_r__36;
      p18_bit_slice_6562 <= p18_data_enable ? p17_bit_slice_6562 : p18_bit_slice_6562;
      p18_bit_slice_6563 <= p18_data_enable ? p17_bit_slice_6563 : p18_bit_slice_6563;
      p18_bit_slice_6564 <= p18_data_enable ? p17_bit_slice_6564 : p18_bit_slice_6564;
      p18_bit_slice_6565 <= p18_data_enable ? p17_bit_slice_6565 : p18_bit_slice_6565;
      p18_bit_slice_6566 <= p18_data_enable ? p17_bit_slice_6566 : p18_bit_slice_6566;
      p18_bit_slice_6567 <= p18_data_enable ? p17_bit_slice_6567 : p18_bit_slice_6567;
      p18_bit_slice_6568 <= p18_data_enable ? p17_bit_slice_6568 : p18_bit_slice_6568;
      p18_bit_slice_6569 <= p18_data_enable ? p17_bit_slice_6569 : p18_bit_slice_6569;
      p18_bit_slice_6570 <= p18_data_enable ? p17_bit_slice_6570 : p18_bit_slice_6570;
      p18_bit_slice_6571 <= p18_data_enable ? p17_bit_slice_6571 : p18_bit_slice_6571;
      p18_bit_slice_6572 <= p18_data_enable ? p17_bit_slice_6572 : p18_bit_slice_6572;
      p18_bit_slice_6573 <= p18_data_enable ? p17_bit_slice_6573 : p18_bit_slice_6573;
      p18_bit_slice_6574 <= p18_data_enable ? p17_bit_slice_6574 : p18_bit_slice_6574;
      p18_bit_slice_6575 <= p18_data_enable ? p17_bit_slice_6575 : p18_bit_slice_6575;
      p19_b <= p19_data_enable ? p18_b : p19_b;
      p19_uge_6652 <= p19_data_enable ? p18_uge_6652 : p19_uge_6652;
      p19_bivisor__1 <= p19_data_enable ? p18_bivisor__1 : p19_bivisor__1;
      p19_uge_6732 <= p19_data_enable ? p18_uge_6732 : p19_uge_6732;
      p19_uge_6810 <= p19_data_enable ? p18_uge_6810 : p19_uge_6810;
      p19_uge_6888 <= p19_data_enable ? p18_uge_6888 : p19_uge_6888;
      p19_uge_6966 <= p19_data_enable ? p18_uge_6966 : p19_uge_6966;
      p19_uge_7044 <= p19_data_enable ? p18_uge_7044 : p19_uge_7044;
      p19_uge_7122 <= p19_data_enable ? p18_uge_7122 : p19_uge_7122;
      p19_uge_7200 <= p19_data_enable ? p18_uge_7200 : p19_uge_7200;
      p19_uge_7278 <= p19_data_enable ? p18_uge_7278 : p19_uge_7278;
      p19_uge_7356 <= p19_data_enable ? p18_uge_7356 : p19_uge_7356;
      p19_uge_7434 <= p19_data_enable ? p18_uge_7434 : p19_uge_7434;
      p19_uge_7512 <= p19_data_enable ? p18_uge_7512 : p19_uge_7512;
      p19_uge_7590 <= p19_data_enable ? p18_uge_7590 : p19_uge_7590;
      p19_uge_7668 <= p19_data_enable ? p18_uge_7668 : p19_uge_7668;
      p19_uge_7746 <= p19_data_enable ? p18_uge_7746 : p19_uge_7746;
      p19_uge_7824 <= p19_data_enable ? p18_uge_7824 : p19_uge_7824;
      p19_uge_7902 <= p19_data_enable ? p18_uge_7902 : p19_uge_7902;
      p19_uge_7980 <= p19_data_enable ? p18_uge_7980 : p19_uge_7980;
      p19_uge_8058 <= p19_data_enable ? uge_8058 : p19_uge_8058;
      p19_r__38 <= p19_data_enable ? r__38 : p19_r__38;
      p19_bit_slice_6563 <= p19_data_enable ? p18_bit_slice_6563 : p19_bit_slice_6563;
      p19_bit_slice_6564 <= p19_data_enable ? p18_bit_slice_6564 : p19_bit_slice_6564;
      p19_bit_slice_6565 <= p19_data_enable ? p18_bit_slice_6565 : p19_bit_slice_6565;
      p19_bit_slice_6566 <= p19_data_enable ? p18_bit_slice_6566 : p19_bit_slice_6566;
      p19_bit_slice_6567 <= p19_data_enable ? p18_bit_slice_6567 : p19_bit_slice_6567;
      p19_bit_slice_6568 <= p19_data_enable ? p18_bit_slice_6568 : p19_bit_slice_6568;
      p19_bit_slice_6569 <= p19_data_enable ? p18_bit_slice_6569 : p19_bit_slice_6569;
      p19_bit_slice_6570 <= p19_data_enable ? p18_bit_slice_6570 : p19_bit_slice_6570;
      p19_bit_slice_6571 <= p19_data_enable ? p18_bit_slice_6571 : p19_bit_slice_6571;
      p19_bit_slice_6572 <= p19_data_enable ? p18_bit_slice_6572 : p19_bit_slice_6572;
      p19_bit_slice_6573 <= p19_data_enable ? p18_bit_slice_6573 : p19_bit_slice_6573;
      p19_bit_slice_6574 <= p19_data_enable ? p18_bit_slice_6574 : p19_bit_slice_6574;
      p19_bit_slice_6575 <= p19_data_enable ? p18_bit_slice_6575 : p19_bit_slice_6575;
      p20_b <= p20_data_enable ? p19_b : p20_b;
      p20_uge_6652 <= p20_data_enable ? p19_uge_6652 : p20_uge_6652;
      p20_bivisor__1 <= p20_data_enable ? p19_bivisor__1 : p20_bivisor__1;
      p20_uge_6732 <= p20_data_enable ? p19_uge_6732 : p20_uge_6732;
      p20_uge_6810 <= p20_data_enable ? p19_uge_6810 : p20_uge_6810;
      p20_uge_6888 <= p20_data_enable ? p19_uge_6888 : p20_uge_6888;
      p20_uge_6966 <= p20_data_enable ? p19_uge_6966 : p20_uge_6966;
      p20_uge_7044 <= p20_data_enable ? p19_uge_7044 : p20_uge_7044;
      p20_uge_7122 <= p20_data_enable ? p19_uge_7122 : p20_uge_7122;
      p20_uge_7200 <= p20_data_enable ? p19_uge_7200 : p20_uge_7200;
      p20_uge_7278 <= p20_data_enable ? p19_uge_7278 : p20_uge_7278;
      p20_uge_7356 <= p20_data_enable ? p19_uge_7356 : p20_uge_7356;
      p20_uge_7434 <= p20_data_enable ? p19_uge_7434 : p20_uge_7434;
      p20_uge_7512 <= p20_data_enable ? p19_uge_7512 : p20_uge_7512;
      p20_uge_7590 <= p20_data_enable ? p19_uge_7590 : p20_uge_7590;
      p20_uge_7668 <= p20_data_enable ? p19_uge_7668 : p20_uge_7668;
      p20_uge_7746 <= p20_data_enable ? p19_uge_7746 : p20_uge_7746;
      p20_uge_7824 <= p20_data_enable ? p19_uge_7824 : p20_uge_7824;
      p20_uge_7902 <= p20_data_enable ? p19_uge_7902 : p20_uge_7902;
      p20_uge_7980 <= p20_data_enable ? p19_uge_7980 : p20_uge_7980;
      p20_uge_8058 <= p20_data_enable ? p19_uge_8058 : p20_uge_8058;
      p20_uge_8136 <= p20_data_enable ? uge_8136 : p20_uge_8136;
      p20_r__40 <= p20_data_enable ? r__40 : p20_r__40;
      p20_bit_slice_6564 <= p20_data_enable ? p19_bit_slice_6564 : p20_bit_slice_6564;
      p20_bit_slice_6565 <= p20_data_enable ? p19_bit_slice_6565 : p20_bit_slice_6565;
      p20_bit_slice_6566 <= p20_data_enable ? p19_bit_slice_6566 : p20_bit_slice_6566;
      p20_bit_slice_6567 <= p20_data_enable ? p19_bit_slice_6567 : p20_bit_slice_6567;
      p20_bit_slice_6568 <= p20_data_enable ? p19_bit_slice_6568 : p20_bit_slice_6568;
      p20_bit_slice_6569 <= p20_data_enable ? p19_bit_slice_6569 : p20_bit_slice_6569;
      p20_bit_slice_6570 <= p20_data_enable ? p19_bit_slice_6570 : p20_bit_slice_6570;
      p20_bit_slice_6571 <= p20_data_enable ? p19_bit_slice_6571 : p20_bit_slice_6571;
      p20_bit_slice_6572 <= p20_data_enable ? p19_bit_slice_6572 : p20_bit_slice_6572;
      p20_bit_slice_6573 <= p20_data_enable ? p19_bit_slice_6573 : p20_bit_slice_6573;
      p20_bit_slice_6574 <= p20_data_enable ? p19_bit_slice_6574 : p20_bit_slice_6574;
      p20_bit_slice_6575 <= p20_data_enable ? p19_bit_slice_6575 : p20_bit_slice_6575;
      p21_b <= p21_data_enable ? p20_b : p21_b;
      p21_uge_6652 <= p21_data_enable ? p20_uge_6652 : p21_uge_6652;
      p21_bivisor__1 <= p21_data_enable ? p20_bivisor__1 : p21_bivisor__1;
      p21_uge_6732 <= p21_data_enable ? p20_uge_6732 : p21_uge_6732;
      p21_uge_6810 <= p21_data_enable ? p20_uge_6810 : p21_uge_6810;
      p21_uge_6888 <= p21_data_enable ? p20_uge_6888 : p21_uge_6888;
      p21_uge_6966 <= p21_data_enable ? p20_uge_6966 : p21_uge_6966;
      p21_uge_7044 <= p21_data_enable ? p20_uge_7044 : p21_uge_7044;
      p21_uge_7122 <= p21_data_enable ? p20_uge_7122 : p21_uge_7122;
      p21_uge_7200 <= p21_data_enable ? p20_uge_7200 : p21_uge_7200;
      p21_uge_7278 <= p21_data_enable ? p20_uge_7278 : p21_uge_7278;
      p21_uge_7356 <= p21_data_enable ? p20_uge_7356 : p21_uge_7356;
      p21_uge_7434 <= p21_data_enable ? p20_uge_7434 : p21_uge_7434;
      p21_uge_7512 <= p21_data_enable ? p20_uge_7512 : p21_uge_7512;
      p21_uge_7590 <= p21_data_enable ? p20_uge_7590 : p21_uge_7590;
      p21_uge_7668 <= p21_data_enable ? p20_uge_7668 : p21_uge_7668;
      p21_uge_7746 <= p21_data_enable ? p20_uge_7746 : p21_uge_7746;
      p21_uge_7824 <= p21_data_enable ? p20_uge_7824 : p21_uge_7824;
      p21_uge_7902 <= p21_data_enable ? p20_uge_7902 : p21_uge_7902;
      p21_uge_7980 <= p21_data_enable ? p20_uge_7980 : p21_uge_7980;
      p21_uge_8058 <= p21_data_enable ? p20_uge_8058 : p21_uge_8058;
      p21_uge_8136 <= p21_data_enable ? p20_uge_8136 : p21_uge_8136;
      p21_uge_8214 <= p21_data_enable ? uge_8214 : p21_uge_8214;
      p21_r__42 <= p21_data_enable ? r__42 : p21_r__42;
      p21_bit_slice_6565 <= p21_data_enable ? p20_bit_slice_6565 : p21_bit_slice_6565;
      p21_bit_slice_6566 <= p21_data_enable ? p20_bit_slice_6566 : p21_bit_slice_6566;
      p21_bit_slice_6567 <= p21_data_enable ? p20_bit_slice_6567 : p21_bit_slice_6567;
      p21_bit_slice_6568 <= p21_data_enable ? p20_bit_slice_6568 : p21_bit_slice_6568;
      p21_bit_slice_6569 <= p21_data_enable ? p20_bit_slice_6569 : p21_bit_slice_6569;
      p21_bit_slice_6570 <= p21_data_enable ? p20_bit_slice_6570 : p21_bit_slice_6570;
      p21_bit_slice_6571 <= p21_data_enable ? p20_bit_slice_6571 : p21_bit_slice_6571;
      p21_bit_slice_6572 <= p21_data_enable ? p20_bit_slice_6572 : p21_bit_slice_6572;
      p21_bit_slice_6573 <= p21_data_enable ? p20_bit_slice_6573 : p21_bit_slice_6573;
      p21_bit_slice_6574 <= p21_data_enable ? p20_bit_slice_6574 : p21_bit_slice_6574;
      p21_bit_slice_6575 <= p21_data_enable ? p20_bit_slice_6575 : p21_bit_slice_6575;
      p22_b <= p22_data_enable ? p21_b : p22_b;
      p22_uge_6652 <= p22_data_enable ? p21_uge_6652 : p22_uge_6652;
      p22_bivisor__1 <= p22_data_enable ? p21_bivisor__1 : p22_bivisor__1;
      p22_uge_6732 <= p22_data_enable ? p21_uge_6732 : p22_uge_6732;
      p22_uge_6810 <= p22_data_enable ? p21_uge_6810 : p22_uge_6810;
      p22_uge_6888 <= p22_data_enable ? p21_uge_6888 : p22_uge_6888;
      p22_uge_6966 <= p22_data_enable ? p21_uge_6966 : p22_uge_6966;
      p22_uge_7044 <= p22_data_enable ? p21_uge_7044 : p22_uge_7044;
      p22_uge_7122 <= p22_data_enable ? p21_uge_7122 : p22_uge_7122;
      p22_uge_7200 <= p22_data_enable ? p21_uge_7200 : p22_uge_7200;
      p22_uge_7278 <= p22_data_enable ? p21_uge_7278 : p22_uge_7278;
      p22_uge_7356 <= p22_data_enable ? p21_uge_7356 : p22_uge_7356;
      p22_uge_7434 <= p22_data_enable ? p21_uge_7434 : p22_uge_7434;
      p22_uge_7512 <= p22_data_enable ? p21_uge_7512 : p22_uge_7512;
      p22_uge_7590 <= p22_data_enable ? p21_uge_7590 : p22_uge_7590;
      p22_uge_7668 <= p22_data_enable ? p21_uge_7668 : p22_uge_7668;
      p22_uge_7746 <= p22_data_enable ? p21_uge_7746 : p22_uge_7746;
      p22_uge_7824 <= p22_data_enable ? p21_uge_7824 : p22_uge_7824;
      p22_uge_7902 <= p22_data_enable ? p21_uge_7902 : p22_uge_7902;
      p22_uge_7980 <= p22_data_enable ? p21_uge_7980 : p22_uge_7980;
      p22_uge_8058 <= p22_data_enable ? p21_uge_8058 : p22_uge_8058;
      p22_uge_8136 <= p22_data_enable ? p21_uge_8136 : p22_uge_8136;
      p22_uge_8214 <= p22_data_enable ? p21_uge_8214 : p22_uge_8214;
      p22_uge_8292 <= p22_data_enable ? uge_8292 : p22_uge_8292;
      p22_r__44 <= p22_data_enable ? r__44 : p22_r__44;
      p22_bit_slice_6566 <= p22_data_enable ? p21_bit_slice_6566 : p22_bit_slice_6566;
      p22_bit_slice_6567 <= p22_data_enable ? p21_bit_slice_6567 : p22_bit_slice_6567;
      p22_bit_slice_6568 <= p22_data_enable ? p21_bit_slice_6568 : p22_bit_slice_6568;
      p22_bit_slice_6569 <= p22_data_enable ? p21_bit_slice_6569 : p22_bit_slice_6569;
      p22_bit_slice_6570 <= p22_data_enable ? p21_bit_slice_6570 : p22_bit_slice_6570;
      p22_bit_slice_6571 <= p22_data_enable ? p21_bit_slice_6571 : p22_bit_slice_6571;
      p22_bit_slice_6572 <= p22_data_enable ? p21_bit_slice_6572 : p22_bit_slice_6572;
      p22_bit_slice_6573 <= p22_data_enable ? p21_bit_slice_6573 : p22_bit_slice_6573;
      p22_bit_slice_6574 <= p22_data_enable ? p21_bit_slice_6574 : p22_bit_slice_6574;
      p22_bit_slice_6575 <= p22_data_enable ? p21_bit_slice_6575 : p22_bit_slice_6575;
      p23_b <= p23_data_enable ? p22_b : p23_b;
      p23_uge_6652 <= p23_data_enable ? p22_uge_6652 : p23_uge_6652;
      p23_bivisor__1 <= p23_data_enable ? p22_bivisor__1 : p23_bivisor__1;
      p23_uge_6732 <= p23_data_enable ? p22_uge_6732 : p23_uge_6732;
      p23_uge_6810 <= p23_data_enable ? p22_uge_6810 : p23_uge_6810;
      p23_uge_6888 <= p23_data_enable ? p22_uge_6888 : p23_uge_6888;
      p23_uge_6966 <= p23_data_enable ? p22_uge_6966 : p23_uge_6966;
      p23_uge_7044 <= p23_data_enable ? p22_uge_7044 : p23_uge_7044;
      p23_uge_7122 <= p23_data_enable ? p22_uge_7122 : p23_uge_7122;
      p23_uge_7200 <= p23_data_enable ? p22_uge_7200 : p23_uge_7200;
      p23_uge_7278 <= p23_data_enable ? p22_uge_7278 : p23_uge_7278;
      p23_uge_7356 <= p23_data_enable ? p22_uge_7356 : p23_uge_7356;
      p23_uge_7434 <= p23_data_enable ? p22_uge_7434 : p23_uge_7434;
      p23_uge_7512 <= p23_data_enable ? p22_uge_7512 : p23_uge_7512;
      p23_uge_7590 <= p23_data_enable ? p22_uge_7590 : p23_uge_7590;
      p23_uge_7668 <= p23_data_enable ? p22_uge_7668 : p23_uge_7668;
      p23_uge_7746 <= p23_data_enable ? p22_uge_7746 : p23_uge_7746;
      p23_uge_7824 <= p23_data_enable ? p22_uge_7824 : p23_uge_7824;
      p23_uge_7902 <= p23_data_enable ? p22_uge_7902 : p23_uge_7902;
      p23_uge_7980 <= p23_data_enable ? p22_uge_7980 : p23_uge_7980;
      p23_uge_8058 <= p23_data_enable ? p22_uge_8058 : p23_uge_8058;
      p23_uge_8136 <= p23_data_enable ? p22_uge_8136 : p23_uge_8136;
      p23_uge_8214 <= p23_data_enable ? p22_uge_8214 : p23_uge_8214;
      p23_uge_8292 <= p23_data_enable ? p22_uge_8292 : p23_uge_8292;
      p23_uge_8370 <= p23_data_enable ? uge_8370 : p23_uge_8370;
      p23_r__46 <= p23_data_enable ? r__46 : p23_r__46;
      p23_bit_slice_6567 <= p23_data_enable ? p22_bit_slice_6567 : p23_bit_slice_6567;
      p23_bit_slice_6568 <= p23_data_enable ? p22_bit_slice_6568 : p23_bit_slice_6568;
      p23_bit_slice_6569 <= p23_data_enable ? p22_bit_slice_6569 : p23_bit_slice_6569;
      p23_bit_slice_6570 <= p23_data_enable ? p22_bit_slice_6570 : p23_bit_slice_6570;
      p23_bit_slice_6571 <= p23_data_enable ? p22_bit_slice_6571 : p23_bit_slice_6571;
      p23_bit_slice_6572 <= p23_data_enable ? p22_bit_slice_6572 : p23_bit_slice_6572;
      p23_bit_slice_6573 <= p23_data_enable ? p22_bit_slice_6573 : p23_bit_slice_6573;
      p23_bit_slice_6574 <= p23_data_enable ? p22_bit_slice_6574 : p23_bit_slice_6574;
      p23_bit_slice_6575 <= p23_data_enable ? p22_bit_slice_6575 : p23_bit_slice_6575;
      p24_b <= p24_data_enable ? p23_b : p24_b;
      p24_uge_6652 <= p24_data_enable ? p23_uge_6652 : p24_uge_6652;
      p24_bivisor__1 <= p24_data_enable ? p23_bivisor__1 : p24_bivisor__1;
      p24_uge_6732 <= p24_data_enable ? p23_uge_6732 : p24_uge_6732;
      p24_uge_6810 <= p24_data_enable ? p23_uge_6810 : p24_uge_6810;
      p24_uge_6888 <= p24_data_enable ? p23_uge_6888 : p24_uge_6888;
      p24_uge_6966 <= p24_data_enable ? p23_uge_6966 : p24_uge_6966;
      p24_uge_7044 <= p24_data_enable ? p23_uge_7044 : p24_uge_7044;
      p24_uge_7122 <= p24_data_enable ? p23_uge_7122 : p24_uge_7122;
      p24_uge_7200 <= p24_data_enable ? p23_uge_7200 : p24_uge_7200;
      p24_uge_7278 <= p24_data_enable ? p23_uge_7278 : p24_uge_7278;
      p24_uge_7356 <= p24_data_enable ? p23_uge_7356 : p24_uge_7356;
      p24_uge_7434 <= p24_data_enable ? p23_uge_7434 : p24_uge_7434;
      p24_uge_7512 <= p24_data_enable ? p23_uge_7512 : p24_uge_7512;
      p24_uge_7590 <= p24_data_enable ? p23_uge_7590 : p24_uge_7590;
      p24_uge_7668 <= p24_data_enable ? p23_uge_7668 : p24_uge_7668;
      p24_uge_7746 <= p24_data_enable ? p23_uge_7746 : p24_uge_7746;
      p24_uge_7824 <= p24_data_enable ? p23_uge_7824 : p24_uge_7824;
      p24_uge_7902 <= p24_data_enable ? p23_uge_7902 : p24_uge_7902;
      p24_uge_7980 <= p24_data_enable ? p23_uge_7980 : p24_uge_7980;
      p24_uge_8058 <= p24_data_enable ? p23_uge_8058 : p24_uge_8058;
      p24_uge_8136 <= p24_data_enable ? p23_uge_8136 : p24_uge_8136;
      p24_uge_8214 <= p24_data_enable ? p23_uge_8214 : p24_uge_8214;
      p24_uge_8292 <= p24_data_enable ? p23_uge_8292 : p24_uge_8292;
      p24_uge_8370 <= p24_data_enable ? p23_uge_8370 : p24_uge_8370;
      p24_uge_8448 <= p24_data_enable ? uge_8448 : p24_uge_8448;
      p24_r__48 <= p24_data_enable ? r__48 : p24_r__48;
      p24_bit_slice_6568 <= p24_data_enable ? p23_bit_slice_6568 : p24_bit_slice_6568;
      p24_bit_slice_6569 <= p24_data_enable ? p23_bit_slice_6569 : p24_bit_slice_6569;
      p24_bit_slice_6570 <= p24_data_enable ? p23_bit_slice_6570 : p24_bit_slice_6570;
      p24_bit_slice_6571 <= p24_data_enable ? p23_bit_slice_6571 : p24_bit_slice_6571;
      p24_bit_slice_6572 <= p24_data_enable ? p23_bit_slice_6572 : p24_bit_slice_6572;
      p24_bit_slice_6573 <= p24_data_enable ? p23_bit_slice_6573 : p24_bit_slice_6573;
      p24_bit_slice_6574 <= p24_data_enable ? p23_bit_slice_6574 : p24_bit_slice_6574;
      p24_bit_slice_6575 <= p24_data_enable ? p23_bit_slice_6575 : p24_bit_slice_6575;
      p25_b <= p25_data_enable ? p24_b : p25_b;
      p25_uge_6652 <= p25_data_enable ? p24_uge_6652 : p25_uge_6652;
      p25_bivisor__1 <= p25_data_enable ? p24_bivisor__1 : p25_bivisor__1;
      p25_uge_6732 <= p25_data_enable ? p24_uge_6732 : p25_uge_6732;
      p25_uge_6810 <= p25_data_enable ? p24_uge_6810 : p25_uge_6810;
      p25_uge_6888 <= p25_data_enable ? p24_uge_6888 : p25_uge_6888;
      p25_uge_6966 <= p25_data_enable ? p24_uge_6966 : p25_uge_6966;
      p25_uge_7044 <= p25_data_enable ? p24_uge_7044 : p25_uge_7044;
      p25_uge_7122 <= p25_data_enable ? p24_uge_7122 : p25_uge_7122;
      p25_uge_7200 <= p25_data_enable ? p24_uge_7200 : p25_uge_7200;
      p25_uge_7278 <= p25_data_enable ? p24_uge_7278 : p25_uge_7278;
      p25_uge_7356 <= p25_data_enable ? p24_uge_7356 : p25_uge_7356;
      p25_uge_7434 <= p25_data_enable ? p24_uge_7434 : p25_uge_7434;
      p25_uge_7512 <= p25_data_enable ? p24_uge_7512 : p25_uge_7512;
      p25_uge_7590 <= p25_data_enable ? p24_uge_7590 : p25_uge_7590;
      p25_uge_7668 <= p25_data_enable ? p24_uge_7668 : p25_uge_7668;
      p25_uge_7746 <= p25_data_enable ? p24_uge_7746 : p25_uge_7746;
      p25_uge_7824 <= p25_data_enable ? p24_uge_7824 : p25_uge_7824;
      p25_uge_7902 <= p25_data_enable ? p24_uge_7902 : p25_uge_7902;
      p25_uge_7980 <= p25_data_enable ? p24_uge_7980 : p25_uge_7980;
      p25_uge_8058 <= p25_data_enable ? p24_uge_8058 : p25_uge_8058;
      p25_uge_8136 <= p25_data_enable ? p24_uge_8136 : p25_uge_8136;
      p25_uge_8214 <= p25_data_enable ? p24_uge_8214 : p25_uge_8214;
      p25_uge_8292 <= p25_data_enable ? p24_uge_8292 : p25_uge_8292;
      p25_uge_8370 <= p25_data_enable ? p24_uge_8370 : p25_uge_8370;
      p25_uge_8448 <= p25_data_enable ? p24_uge_8448 : p25_uge_8448;
      p25_uge_8526 <= p25_data_enable ? uge_8526 : p25_uge_8526;
      p25_r__50 <= p25_data_enable ? r__50 : p25_r__50;
      p25_bit_slice_6569 <= p25_data_enable ? p24_bit_slice_6569 : p25_bit_slice_6569;
      p25_bit_slice_6570 <= p25_data_enable ? p24_bit_slice_6570 : p25_bit_slice_6570;
      p25_bit_slice_6571 <= p25_data_enable ? p24_bit_slice_6571 : p25_bit_slice_6571;
      p25_bit_slice_6572 <= p25_data_enable ? p24_bit_slice_6572 : p25_bit_slice_6572;
      p25_bit_slice_6573 <= p25_data_enable ? p24_bit_slice_6573 : p25_bit_slice_6573;
      p25_bit_slice_6574 <= p25_data_enable ? p24_bit_slice_6574 : p25_bit_slice_6574;
      p25_bit_slice_6575 <= p25_data_enable ? p24_bit_slice_6575 : p25_bit_slice_6575;
      p26_b <= p26_data_enable ? p25_b : p26_b;
      p26_uge_6652 <= p26_data_enable ? p25_uge_6652 : p26_uge_6652;
      p26_bivisor__1 <= p26_data_enable ? p25_bivisor__1 : p26_bivisor__1;
      p26_uge_6732 <= p26_data_enable ? p25_uge_6732 : p26_uge_6732;
      p26_uge_6810 <= p26_data_enable ? p25_uge_6810 : p26_uge_6810;
      p26_uge_6888 <= p26_data_enable ? p25_uge_6888 : p26_uge_6888;
      p26_uge_6966 <= p26_data_enable ? p25_uge_6966 : p26_uge_6966;
      p26_uge_7044 <= p26_data_enable ? p25_uge_7044 : p26_uge_7044;
      p26_uge_7122 <= p26_data_enable ? p25_uge_7122 : p26_uge_7122;
      p26_uge_7200 <= p26_data_enable ? p25_uge_7200 : p26_uge_7200;
      p26_uge_7278 <= p26_data_enable ? p25_uge_7278 : p26_uge_7278;
      p26_uge_7356 <= p26_data_enable ? p25_uge_7356 : p26_uge_7356;
      p26_uge_7434 <= p26_data_enable ? p25_uge_7434 : p26_uge_7434;
      p26_uge_7512 <= p26_data_enable ? p25_uge_7512 : p26_uge_7512;
      p26_uge_7590 <= p26_data_enable ? p25_uge_7590 : p26_uge_7590;
      p26_uge_7668 <= p26_data_enable ? p25_uge_7668 : p26_uge_7668;
      p26_uge_7746 <= p26_data_enable ? p25_uge_7746 : p26_uge_7746;
      p26_uge_7824 <= p26_data_enable ? p25_uge_7824 : p26_uge_7824;
      p26_uge_7902 <= p26_data_enable ? p25_uge_7902 : p26_uge_7902;
      p26_uge_7980 <= p26_data_enable ? p25_uge_7980 : p26_uge_7980;
      p26_uge_8058 <= p26_data_enable ? p25_uge_8058 : p26_uge_8058;
      p26_uge_8136 <= p26_data_enable ? p25_uge_8136 : p26_uge_8136;
      p26_uge_8214 <= p26_data_enable ? p25_uge_8214 : p26_uge_8214;
      p26_uge_8292 <= p26_data_enable ? p25_uge_8292 : p26_uge_8292;
      p26_uge_8370 <= p26_data_enable ? p25_uge_8370 : p26_uge_8370;
      p26_uge_8448 <= p26_data_enable ? p25_uge_8448 : p26_uge_8448;
      p26_uge_8526 <= p26_data_enable ? p25_uge_8526 : p26_uge_8526;
      p26_uge_8604 <= p26_data_enable ? uge_8604 : p26_uge_8604;
      p26_r__52 <= p26_data_enable ? r__52 : p26_r__52;
      p26_bit_slice_6570 <= p26_data_enable ? p25_bit_slice_6570 : p26_bit_slice_6570;
      p26_bit_slice_6571 <= p26_data_enable ? p25_bit_slice_6571 : p26_bit_slice_6571;
      p26_bit_slice_6572 <= p26_data_enable ? p25_bit_slice_6572 : p26_bit_slice_6572;
      p26_bit_slice_6573 <= p26_data_enable ? p25_bit_slice_6573 : p26_bit_slice_6573;
      p26_bit_slice_6574 <= p26_data_enable ? p25_bit_slice_6574 : p26_bit_slice_6574;
      p26_bit_slice_6575 <= p26_data_enable ? p25_bit_slice_6575 : p26_bit_slice_6575;
      p27_b <= p27_data_enable ? p26_b : p27_b;
      p27_uge_6652 <= p27_data_enable ? p26_uge_6652 : p27_uge_6652;
      p27_bivisor__1 <= p27_data_enable ? p26_bivisor__1 : p27_bivisor__1;
      p27_uge_6732 <= p27_data_enable ? p26_uge_6732 : p27_uge_6732;
      p27_uge_6810 <= p27_data_enable ? p26_uge_6810 : p27_uge_6810;
      p27_uge_6888 <= p27_data_enable ? p26_uge_6888 : p27_uge_6888;
      p27_uge_6966 <= p27_data_enable ? p26_uge_6966 : p27_uge_6966;
      p27_uge_7044 <= p27_data_enable ? p26_uge_7044 : p27_uge_7044;
      p27_uge_7122 <= p27_data_enable ? p26_uge_7122 : p27_uge_7122;
      p27_uge_7200 <= p27_data_enable ? p26_uge_7200 : p27_uge_7200;
      p27_uge_7278 <= p27_data_enable ? p26_uge_7278 : p27_uge_7278;
      p27_uge_7356 <= p27_data_enable ? p26_uge_7356 : p27_uge_7356;
      p27_uge_7434 <= p27_data_enable ? p26_uge_7434 : p27_uge_7434;
      p27_uge_7512 <= p27_data_enable ? p26_uge_7512 : p27_uge_7512;
      p27_uge_7590 <= p27_data_enable ? p26_uge_7590 : p27_uge_7590;
      p27_uge_7668 <= p27_data_enable ? p26_uge_7668 : p27_uge_7668;
      p27_uge_7746 <= p27_data_enable ? p26_uge_7746 : p27_uge_7746;
      p27_uge_7824 <= p27_data_enable ? p26_uge_7824 : p27_uge_7824;
      p27_uge_7902 <= p27_data_enable ? p26_uge_7902 : p27_uge_7902;
      p27_uge_7980 <= p27_data_enable ? p26_uge_7980 : p27_uge_7980;
      p27_uge_8058 <= p27_data_enable ? p26_uge_8058 : p27_uge_8058;
      p27_uge_8136 <= p27_data_enable ? p26_uge_8136 : p27_uge_8136;
      p27_uge_8214 <= p27_data_enable ? p26_uge_8214 : p27_uge_8214;
      p27_uge_8292 <= p27_data_enable ? p26_uge_8292 : p27_uge_8292;
      p27_uge_8370 <= p27_data_enable ? p26_uge_8370 : p27_uge_8370;
      p27_uge_8448 <= p27_data_enable ? p26_uge_8448 : p27_uge_8448;
      p27_uge_8526 <= p27_data_enable ? p26_uge_8526 : p27_uge_8526;
      p27_uge_8604 <= p27_data_enable ? p26_uge_8604 : p27_uge_8604;
      p27_uge_8682 <= p27_data_enable ? uge_8682 : p27_uge_8682;
      p27_r__54 <= p27_data_enable ? r__54 : p27_r__54;
      p27_bit_slice_6571 <= p27_data_enable ? p26_bit_slice_6571 : p27_bit_slice_6571;
      p27_bit_slice_6572 <= p27_data_enable ? p26_bit_slice_6572 : p27_bit_slice_6572;
      p27_bit_slice_6573 <= p27_data_enable ? p26_bit_slice_6573 : p27_bit_slice_6573;
      p27_bit_slice_6574 <= p27_data_enable ? p26_bit_slice_6574 : p27_bit_slice_6574;
      p27_bit_slice_6575 <= p27_data_enable ? p26_bit_slice_6575 : p27_bit_slice_6575;
      p28_b <= p28_data_enable ? p27_b : p28_b;
      p28_uge_6652 <= p28_data_enable ? p27_uge_6652 : p28_uge_6652;
      p28_bivisor__1 <= p28_data_enable ? p27_bivisor__1 : p28_bivisor__1;
      p28_uge_6732 <= p28_data_enable ? p27_uge_6732 : p28_uge_6732;
      p28_uge_6810 <= p28_data_enable ? p27_uge_6810 : p28_uge_6810;
      p28_uge_6888 <= p28_data_enable ? p27_uge_6888 : p28_uge_6888;
      p28_uge_6966 <= p28_data_enable ? p27_uge_6966 : p28_uge_6966;
      p28_uge_7044 <= p28_data_enable ? p27_uge_7044 : p28_uge_7044;
      p28_uge_7122 <= p28_data_enable ? p27_uge_7122 : p28_uge_7122;
      p28_uge_7200 <= p28_data_enable ? p27_uge_7200 : p28_uge_7200;
      p28_uge_7278 <= p28_data_enable ? p27_uge_7278 : p28_uge_7278;
      p28_uge_7356 <= p28_data_enable ? p27_uge_7356 : p28_uge_7356;
      p28_uge_7434 <= p28_data_enable ? p27_uge_7434 : p28_uge_7434;
      p28_uge_7512 <= p28_data_enable ? p27_uge_7512 : p28_uge_7512;
      p28_uge_7590 <= p28_data_enable ? p27_uge_7590 : p28_uge_7590;
      p28_uge_7668 <= p28_data_enable ? p27_uge_7668 : p28_uge_7668;
      p28_uge_7746 <= p28_data_enable ? p27_uge_7746 : p28_uge_7746;
      p28_uge_7824 <= p28_data_enable ? p27_uge_7824 : p28_uge_7824;
      p28_uge_7902 <= p28_data_enable ? p27_uge_7902 : p28_uge_7902;
      p28_uge_7980 <= p28_data_enable ? p27_uge_7980 : p28_uge_7980;
      p28_uge_8058 <= p28_data_enable ? p27_uge_8058 : p28_uge_8058;
      p28_uge_8136 <= p28_data_enable ? p27_uge_8136 : p28_uge_8136;
      p28_uge_8214 <= p28_data_enable ? p27_uge_8214 : p28_uge_8214;
      p28_uge_8292 <= p28_data_enable ? p27_uge_8292 : p28_uge_8292;
      p28_uge_8370 <= p28_data_enable ? p27_uge_8370 : p28_uge_8370;
      p28_uge_8448 <= p28_data_enable ? p27_uge_8448 : p28_uge_8448;
      p28_uge_8526 <= p28_data_enable ? p27_uge_8526 : p28_uge_8526;
      p28_uge_8604 <= p28_data_enable ? p27_uge_8604 : p28_uge_8604;
      p28_uge_8682 <= p28_data_enable ? p27_uge_8682 : p28_uge_8682;
      p28_uge_8760 <= p28_data_enable ? uge_8760 : p28_uge_8760;
      p28_r__56 <= p28_data_enable ? r__56 : p28_r__56;
      p28_bit_slice_6572 <= p28_data_enable ? p27_bit_slice_6572 : p28_bit_slice_6572;
      p28_bit_slice_6573 <= p28_data_enable ? p27_bit_slice_6573 : p28_bit_slice_6573;
      p28_bit_slice_6574 <= p28_data_enable ? p27_bit_slice_6574 : p28_bit_slice_6574;
      p28_bit_slice_6575 <= p28_data_enable ? p27_bit_slice_6575 : p28_bit_slice_6575;
      p29_b <= p29_data_enable ? p28_b : p29_b;
      p29_uge_6652 <= p29_data_enable ? p28_uge_6652 : p29_uge_6652;
      p29_bivisor__1 <= p29_data_enable ? p28_bivisor__1 : p29_bivisor__1;
      p29_uge_6732 <= p29_data_enable ? p28_uge_6732 : p29_uge_6732;
      p29_uge_6810 <= p29_data_enable ? p28_uge_6810 : p29_uge_6810;
      p29_uge_6888 <= p29_data_enable ? p28_uge_6888 : p29_uge_6888;
      p29_uge_6966 <= p29_data_enable ? p28_uge_6966 : p29_uge_6966;
      p29_uge_7044 <= p29_data_enable ? p28_uge_7044 : p29_uge_7044;
      p29_uge_7122 <= p29_data_enable ? p28_uge_7122 : p29_uge_7122;
      p29_uge_7200 <= p29_data_enable ? p28_uge_7200 : p29_uge_7200;
      p29_uge_7278 <= p29_data_enable ? p28_uge_7278 : p29_uge_7278;
      p29_uge_7356 <= p29_data_enable ? p28_uge_7356 : p29_uge_7356;
      p29_uge_7434 <= p29_data_enable ? p28_uge_7434 : p29_uge_7434;
      p29_uge_7512 <= p29_data_enable ? p28_uge_7512 : p29_uge_7512;
      p29_uge_7590 <= p29_data_enable ? p28_uge_7590 : p29_uge_7590;
      p29_uge_7668 <= p29_data_enable ? p28_uge_7668 : p29_uge_7668;
      p29_uge_7746 <= p29_data_enable ? p28_uge_7746 : p29_uge_7746;
      p29_uge_7824 <= p29_data_enable ? p28_uge_7824 : p29_uge_7824;
      p29_uge_7902 <= p29_data_enable ? p28_uge_7902 : p29_uge_7902;
      p29_uge_7980 <= p29_data_enable ? p28_uge_7980 : p29_uge_7980;
      p29_uge_8058 <= p29_data_enable ? p28_uge_8058 : p29_uge_8058;
      p29_uge_8136 <= p29_data_enable ? p28_uge_8136 : p29_uge_8136;
      p29_uge_8214 <= p29_data_enable ? p28_uge_8214 : p29_uge_8214;
      p29_uge_8292 <= p29_data_enable ? p28_uge_8292 : p29_uge_8292;
      p29_uge_8370 <= p29_data_enable ? p28_uge_8370 : p29_uge_8370;
      p29_uge_8448 <= p29_data_enable ? p28_uge_8448 : p29_uge_8448;
      p29_uge_8526 <= p29_data_enable ? p28_uge_8526 : p29_uge_8526;
      p29_uge_8604 <= p29_data_enable ? p28_uge_8604 : p29_uge_8604;
      p29_uge_8682 <= p29_data_enable ? p28_uge_8682 : p29_uge_8682;
      p29_uge_8760 <= p29_data_enable ? p28_uge_8760 : p29_uge_8760;
      p29_uge_8838 <= p29_data_enable ? uge_8838 : p29_uge_8838;
      p29_r__58 <= p29_data_enable ? r__58 : p29_r__58;
      p29_bit_slice_6573 <= p29_data_enable ? p28_bit_slice_6573 : p29_bit_slice_6573;
      p29_bit_slice_6574 <= p29_data_enable ? p28_bit_slice_6574 : p29_bit_slice_6574;
      p29_bit_slice_6575 <= p29_data_enable ? p28_bit_slice_6575 : p29_bit_slice_6575;
      p30_b <= p30_data_enable ? p29_b : p30_b;
      p30_uge_6652 <= p30_data_enable ? p29_uge_6652 : p30_uge_6652;
      p30_bivisor__1 <= p30_data_enable ? p29_bivisor__1 : p30_bivisor__1;
      p30_uge_6732 <= p30_data_enable ? p29_uge_6732 : p30_uge_6732;
      p30_uge_6810 <= p30_data_enable ? p29_uge_6810 : p30_uge_6810;
      p30_uge_6888 <= p30_data_enable ? p29_uge_6888 : p30_uge_6888;
      p30_uge_6966 <= p30_data_enable ? p29_uge_6966 : p30_uge_6966;
      p30_uge_7044 <= p30_data_enable ? p29_uge_7044 : p30_uge_7044;
      p30_uge_7122 <= p30_data_enable ? p29_uge_7122 : p30_uge_7122;
      p30_uge_7200 <= p30_data_enable ? p29_uge_7200 : p30_uge_7200;
      p30_uge_7278 <= p30_data_enable ? p29_uge_7278 : p30_uge_7278;
      p30_uge_7356 <= p30_data_enable ? p29_uge_7356 : p30_uge_7356;
      p30_uge_7434 <= p30_data_enable ? p29_uge_7434 : p30_uge_7434;
      p30_uge_7512 <= p30_data_enable ? p29_uge_7512 : p30_uge_7512;
      p30_uge_7590 <= p30_data_enable ? p29_uge_7590 : p30_uge_7590;
      p30_uge_7668 <= p30_data_enable ? p29_uge_7668 : p30_uge_7668;
      p30_uge_7746 <= p30_data_enable ? p29_uge_7746 : p30_uge_7746;
      p30_uge_7824 <= p30_data_enable ? p29_uge_7824 : p30_uge_7824;
      p30_uge_7902 <= p30_data_enable ? p29_uge_7902 : p30_uge_7902;
      p30_uge_7980 <= p30_data_enable ? p29_uge_7980 : p30_uge_7980;
      p30_uge_8058 <= p30_data_enable ? p29_uge_8058 : p30_uge_8058;
      p30_uge_8136 <= p30_data_enable ? p29_uge_8136 : p30_uge_8136;
      p30_uge_8214 <= p30_data_enable ? p29_uge_8214 : p30_uge_8214;
      p30_uge_8292 <= p30_data_enable ? p29_uge_8292 : p30_uge_8292;
      p30_uge_8370 <= p30_data_enable ? p29_uge_8370 : p30_uge_8370;
      p30_uge_8448 <= p30_data_enable ? p29_uge_8448 : p30_uge_8448;
      p30_uge_8526 <= p30_data_enable ? p29_uge_8526 : p30_uge_8526;
      p30_uge_8604 <= p30_data_enable ? p29_uge_8604 : p30_uge_8604;
      p30_uge_8682 <= p30_data_enable ? p29_uge_8682 : p30_uge_8682;
      p30_uge_8760 <= p30_data_enable ? p29_uge_8760 : p30_uge_8760;
      p30_uge_8838 <= p30_data_enable ? p29_uge_8838 : p30_uge_8838;
      p30_uge_8916 <= p30_data_enable ? uge_8916 : p30_uge_8916;
      p30_r__60 <= p30_data_enable ? r__60 : p30_r__60;
      p30_bit_slice_6574 <= p30_data_enable ? p29_bit_slice_6574 : p30_bit_slice_6574;
      p30_bit_slice_6575 <= p30_data_enable ? p29_bit_slice_6575 : p30_bit_slice_6575;
      p31_uge_6652 <= p31_data_enable ? p30_uge_6652 : p31_uge_6652;
      p31_bivisor__1 <= p31_data_enable ? p30_bivisor__1 : p31_bivisor__1;
      p31_uge_6732 <= p31_data_enable ? p30_uge_6732 : p31_uge_6732;
      p31_uge_6810 <= p31_data_enable ? p30_uge_6810 : p31_uge_6810;
      p31_uge_6888 <= p31_data_enable ? p30_uge_6888 : p31_uge_6888;
      p31_uge_6966 <= p31_data_enable ? p30_uge_6966 : p31_uge_6966;
      p31_uge_7044 <= p31_data_enable ? p30_uge_7044 : p31_uge_7044;
      p31_uge_7122 <= p31_data_enable ? p30_uge_7122 : p31_uge_7122;
      p31_uge_7200 <= p31_data_enable ? p30_uge_7200 : p31_uge_7200;
      p31_uge_7278 <= p31_data_enable ? p30_uge_7278 : p31_uge_7278;
      p31_uge_7356 <= p31_data_enable ? p30_uge_7356 : p31_uge_7356;
      p31_uge_7434 <= p31_data_enable ? p30_uge_7434 : p31_uge_7434;
      p31_uge_7512 <= p31_data_enable ? p30_uge_7512 : p31_uge_7512;
      p31_uge_7590 <= p31_data_enable ? p30_uge_7590 : p31_uge_7590;
      p31_uge_7668 <= p31_data_enable ? p30_uge_7668 : p31_uge_7668;
      p31_uge_7746 <= p31_data_enable ? p30_uge_7746 : p31_uge_7746;
      p31_uge_7824 <= p31_data_enable ? p30_uge_7824 : p31_uge_7824;
      p31_uge_7902 <= p31_data_enable ? p30_uge_7902 : p31_uge_7902;
      p31_uge_7980 <= p31_data_enable ? p30_uge_7980 : p31_uge_7980;
      p31_uge_8058 <= p31_data_enable ? p30_uge_8058 : p31_uge_8058;
      p31_uge_8136 <= p31_data_enable ? p30_uge_8136 : p31_uge_8136;
      p31_uge_8214 <= p31_data_enable ? p30_uge_8214 : p31_uge_8214;
      p31_uge_8292 <= p31_data_enable ? p30_uge_8292 : p31_uge_8292;
      p31_uge_8370 <= p31_data_enable ? p30_uge_8370 : p31_uge_8370;
      p31_uge_8448 <= p31_data_enable ? p30_uge_8448 : p31_uge_8448;
      p31_uge_8526 <= p31_data_enable ? p30_uge_8526 : p31_uge_8526;
      p31_uge_8604 <= p31_data_enable ? p30_uge_8604 : p31_uge_8604;
      p31_uge_8682 <= p31_data_enable ? p30_uge_8682 : p31_uge_8682;
      p31_uge_8760 <= p31_data_enable ? p30_uge_8760 : p31_uge_8760;
      p31_uge_8838 <= p31_data_enable ? p30_uge_8838 : p31_uge_8838;
      p31_uge_8916 <= p31_data_enable ? p30_uge_8916 : p31_uge_8916;
      p31_uge_8994 <= p31_data_enable ? uge_8994 : p31_uge_8994;
      p31_r__62 <= p31_data_enable ? r__62 : p31_r__62;
      p31_bit_slice_6575 <= p31_data_enable ? p30_bit_slice_6575 : p31_bit_slice_6575;
      p0_valid <= p0_enable ? xls_float_ips__lhs_vld : p0_valid;
      p1_valid <= p1_enable ? p1_stage_done : p1_valid;
      p2_valid <= p2_enable ? p1_valid : p2_valid;
      p3_valid <= p3_enable ? p2_valid : p3_valid;
      p4_valid <= p4_enable ? p3_valid : p4_valid;
      p5_valid <= p5_enable ? p4_valid : p5_valid;
      p6_valid <= p6_enable ? p5_valid : p6_valid;
      p7_valid <= p7_enable ? p6_valid : p7_valid;
      p8_valid <= p8_enable ? p7_valid : p8_valid;
      p9_valid <= p9_enable ? p8_valid : p9_valid;
      p10_valid <= p10_enable ? p9_valid : p10_valid;
      p11_valid <= p11_enable ? p10_valid : p11_valid;
      p12_valid <= p12_enable ? p11_valid : p12_valid;
      p13_valid <= p13_enable ? p12_valid : p13_valid;
      p14_valid <= p14_enable ? p13_valid : p14_valid;
      p15_valid <= p15_enable ? p14_valid : p15_valid;
      p16_valid <= p16_enable ? p15_valid : p16_valid;
      p17_valid <= p17_enable ? p16_valid : p17_valid;
      p18_valid <= p18_enable ? p17_valid : p18_valid;
      p19_valid <= p19_enable ? p18_valid : p19_valid;
      p20_valid <= p20_enable ? p19_valid : p20_valid;
      p21_valid <= p21_enable ? p20_valid : p21_valid;
      p22_valid <= p22_enable ? p21_valid : p22_valid;
      p23_valid <= p23_enable ? p22_valid : p23_valid;
      p24_valid <= p24_enable ? p23_valid : p24_valid;
      p25_valid <= p25_enable ? p24_valid : p25_valid;
      p26_valid <= p26_enable ? p25_valid : p26_valid;
      p27_valid <= p27_enable ? p26_valid : p27_valid;
      p28_valid <= p28_enable ? p27_valid : p28_valid;
      p29_valid <= p29_enable ? p28_valid : p29_valid;
      p30_valid <= p30_enable ? p29_valid : p30_valid;
      p31_valid <= p31_enable ? p30_valid : p31_valid;
      p32_valid <= p32_enable ? p32_stage_done : p32_valid;
      p33_valid <= p33_enable ? p32_valid : p33_valid;
      p34_valid <= p34_enable ? p33_valid : p34_valid;
      __xls_float_ips__result_reg <= xls_float_ips__result_load_en ? q__32 : __xls_float_ips__result_reg;
      __xls_float_ips__result_valid_reg <= xls_float_ips__result_valid_load_en ? p31_valid : __xls_float_ips__result_valid_reg;
    end
  end
  assign xls_float_ips__result = __xls_float_ips__result_reg;
  assign xls_float_ips__result_vld = __xls_float_ips__result_valid_reg;
  assign xls_float_ips__lhs_rdy = p0_data_enable;
  assign xls_float_ips__rhs_rdy = p1_data_enable;
endmodule
module __xls_float_ips__extf_0_next(
  input wire clk,
  input wire rst,
  input wire [31:0] xls_float_ips__ins,
  input wire xls_float_ips__ins_vld,
  input wire xls_float_ips__outs_rdy,
  output wire [63:0] xls_float_ips__outs,
  output wire xls_float_ips__outs_vld,
  output wire xls_float_ips__ins_rdy
);
  function automatic priority_sel_1b_2way (input reg [1:0] sel, input reg case0, input reg case1, input reg default_value);
    begin
      casez (sel)
        2'b?1: begin
          priority_sel_1b_2way = case0;
        end
        2'b10: begin
          priority_sel_1b_2way = case1;
        end
        2'b00: begin
          priority_sel_1b_2way = default_value;
        end
        default: begin
          // Propagate X
          priority_sel_1b_2way = 1'dx;
        end
      endcase
    end
  endfunction
  function automatic [10:0] priority_sel_11b_2way (input reg [1:0] sel, input reg [10:0] case0, input reg [10:0] case1, input reg [10:0] default_value);
    begin
      casez (sel)
        2'b?1: begin
          priority_sel_11b_2way = case0;
        end
        2'b10: begin
          priority_sel_11b_2way = case1;
        end
        2'b00: begin
          priority_sel_11b_2way = default_value;
        end
        default: begin
          // Propagate X
          priority_sel_11b_2way = 11'dx;
        end
      endcase
    end
  endfunction
  wire [63:0] __xls_float_ips__outs_reg_init = {1'h0, 11'h000, 52'h0_0000_0000_0000};
  reg [63:0] __xls_float_ips__outs_reg;
  reg __xls_float_ips__outs_valid_reg;
  wire [7:0] a_bexp__1;
  wire eq_830;
  wire [22:0] a_fraction__1;
  wire [7:0] EXPR_MASK;
  wire eq_836;
  wire eq_837;
  wire [8:0] arom_exp;
  wire nor_846;
  wire xls_float_ips__outs_valid_inv;
  wire a_sign;
  wire [10:0] TO_EXP_OFFSET;
  wire xls_float_ips__outs_valid_load_en;
  wire [10:0] to_bexp;
  wire xls_float_ips__outs_load_en;
  wire [51:0] concat_867;
  wire p0_stage_done;
  wire [63:0] __xls_float_ips__outs_buf;
  assign a_bexp__1 = xls_float_ips__ins[30:23];
  assign eq_830 = a_bexp__1 == 8'h00;
  assign a_fraction__1 = xls_float_ips__ins[22:0];
  assign EXPR_MASK = 8'hff;
  assign eq_836 = a_fraction__1 == 23'h00_0000;
  assign eq_837 = a_bexp__1 == EXPR_MASK;
  assign arom_exp = {1'h0, a_bexp__1} + 9'h181;
  assign nor_846 = ~(~eq_837 | eq_836);
  assign xls_float_ips__outs_valid_inv = ~__xls_float_ips__outs_valid_reg;
  assign a_sign = xls_float_ips__ins[31:31];
  assign TO_EXP_OFFSET = 11'h3ff;
  assign xls_float_ips__outs_valid_load_en = xls_float_ips__outs_rdy | xls_float_ips__outs_valid_inv;
  assign to_bexp = {{2{arom_exp[8]}}, arom_exp} + TO_EXP_OFFSET;
  assign xls_float_ips__outs_load_en = xls_float_ips__ins_vld & xls_float_ips__outs_valid_load_en;
  assign concat_867 = {priority_sel_1b_2way({~(~eq_830 | eq_836) | eq_830 & eq_836 | eq_837 & eq_836, nor_846}, 1'h1, 1'h0, a_fraction__1[22]), a_fraction__1[21:0] & {22{~(eq_837 | eq_830)}}, 29'h0000_0000};
  assign p0_stage_done = xls_float_ips__ins_vld & xls_float_ips__outs_load_en;
  assign __xls_float_ips__outs_buf = {~(nor_846 | ~a_sign), priority_sel_11b_2way({eq_830, eq_837}, 11'h7ff, 11'h000, to_bexp), concat_867};
  always @ (posedge clk) begin
    if (rst) begin
      __xls_float_ips__outs_reg <= __xls_float_ips__outs_reg_init;
      __xls_float_ips__outs_valid_reg <= 1'h0;
    end else begin
      __xls_float_ips__outs_reg <= xls_float_ips__outs_load_en ? __xls_float_ips__outs_buf : __xls_float_ips__outs_reg;
      __xls_float_ips__outs_valid_reg <= xls_float_ips__outs_valid_load_en ? xls_float_ips__ins_vld : __xls_float_ips__outs_valid_reg;
    end
  end
  assign xls_float_ips__outs = __xls_float_ips__outs_reg;
  assign xls_float_ips__outs_vld = __xls_float_ips__outs_valid_reg;
  assign xls_float_ips__ins_rdy = p0_stage_done;
endmodule
module __xls_float_ips__fptosi_0_next(
  input wire clk,
  input wire rst,
  input wire [31:0] xls_float_ips__ins,
  input wire xls_float_ips__ins_vld,
  input wire xls_float_ips__outs_rdy,
  output wire [31:0] xls_float_ips__outs,
  output wire xls_float_ips__outs_vld,
  output wire xls_float_ips__ins_rdy
);
  reg [7:0] p0_a_bexp__2;
  reg [22:0] p0_a_fraction__2;
  reg p0_a_sign__1;
  reg [22:0] p1_a_fraction__2;
  reg [8:0] p1_add_583;
  reg p1_or_594;
  reg p1_eq_597;
  reg p1_a_sign__1;
  reg p1_or_600;
  reg p2_eq_597;
  reg [31:0] p2_sel_625;
  reg p2_not_626;
  reg p2_a_sign__1;
  reg p2_or_600;
  reg p3_a_sign__1;
  reg [31:0] p3_result;
  reg p0_valid;
  reg p1_valid;
  reg p2_valid;
  reg p3_valid;
  reg [31:0] __xls_float_ips__outs_reg;
  reg __xls_float_ips__outs_valid_reg;
  wire xls_float_ips__outs_valid_inv;
  wire xls_float_ips__outs_valid_load_en;
  wire xls_float_ips__outs_load_en;
  wire p4_stage_done;
  wire p4_not_valid;
  wire p3_enable;
  wire p3_data_enable;
  wire p3_not_valid;
  wire p2_enable;
  wire p2_data_enable;
  wire p2_not_valid;
  wire [31:0] fraction;
  wire [31:0] effective_exp;
  wire [7:0] uexp;
  wire [7:0] subnormal_exp;
  wire eq_588;
  wire p1_enable;
  wire [31:0] INT_MAX;
  wire [31:0] INT_MIN;
  wire ne_589;
  wire [7:0] exp;
  wire p1_data_enable;
  wire p1_not_valid;
  wire exp_oob;
  wire p0_enable;
  wire [31:0] result;
  wire [31:0] sel_625;
  wire not_626;
  wire [8:0] add_583;
  wire or_594;
  wire eq_597;
  wire or_600;
  wire [7:0] a_bexp__2;
  wire p0_data_enable;
  wire [22:0] a_fraction__2;
  wire a_sign__1;
  wire [31:0] result__2;
  assign xls_float_ips__outs_valid_inv = ~__xls_float_ips__outs_valid_reg;
  assign xls_float_ips__outs_valid_load_en = xls_float_ips__outs_rdy | xls_float_ips__outs_valid_inv;
  assign xls_float_ips__outs_load_en = p3_valid & xls_float_ips__outs_valid_load_en;
  assign p4_stage_done = p3_valid & xls_float_ips__outs_load_en;
  assign p4_not_valid = ~p3_valid;
  assign p3_enable = p4_stage_done | p4_not_valid;
  assign p3_data_enable = p3_enable & p2_valid;
  assign p3_not_valid = ~p2_valid;
  assign p2_enable = p3_data_enable | p3_not_valid;
  assign p2_data_enable = p2_enable & p1_valid;
  assign p2_not_valid = ~p1_valid;
  assign fraction = {9'h001, p1_a_fraction__2};
  assign effective_exp = {{23{p1_add_583[8]}}, p1_add_583};
  assign uexp = p0_a_bexp__2 + 8'h81;
  assign subnormal_exp = 8'h82;
  assign eq_588 = p0_a_bexp__2 == 8'hff;
  assign p1_enable = p2_data_enable | p2_not_valid;
  assign INT_MAX = 32'h7fff_ffff;
  assign INT_MIN = 32'h8000_0000;
  assign ne_589 = p0_a_fraction__2 != 23'h00_0000;
  assign exp = p0_a_bexp__2 == 8'h00 ? subnormal_exp : uexp;
  assign p1_data_enable = p1_enable & p0_valid;
  assign p1_not_valid = ~p0_valid;
  assign exp_oob = $signed(exp) >= $signed(8'h1f);
  assign p0_enable = p1_data_enable | p1_not_valid;
  assign result = p2_or_600 ? (p2_a_sign__1 ? INT_MIN : INT_MAX) : (p2_eq_597 ? 32'h0000_0001 : p2_sel_625) & {32{p2_not_626}};
  assign sel_625 = effective_exp[31] ? (-effective_exp >= 32'h0000_0020 ? 32'h0000_0000 : fraction >> -effective_exp) : ($signed(p1_add_583) > $signed(9'h000) ? (effective_exp >= 32'h0000_0020 ? 32'h0000_0000 : fraction << effective_exp) : fraction);
  assign not_626 = ~p1_or_594;
  assign add_583 = {{1{uexp[7]}}, uexp} + 9'h1e9;
  assign or_594 = eq_588 & ne_589 | exp[7];
  assign eq_597 = p0_a_bexp__2 == 8'h7f;
  assign or_600 = exp_oob | ~(~eq_588 | ne_589);
  assign a_bexp__2 = xls_float_ips__ins[30:23];
  assign p0_data_enable = p0_enable & xls_float_ips__ins_vld;
  assign a_fraction__2 = xls_float_ips__ins[22:0];
  assign a_sign__1 = xls_float_ips__ins[31:31];
  assign result__2 = p3_a_sign__1 ? -p3_result : p3_result;
  always @ (posedge clk) begin
    if (rst) begin
      p0_a_bexp__2 <= 8'h00;
      p0_a_fraction__2 <= 23'h00_0000;
      p0_a_sign__1 <= 1'h0;
      p1_a_fraction__2 <= 23'h00_0000;
      p1_add_583 <= 9'h000;
      p1_or_594 <= 1'h0;
      p1_eq_597 <= 1'h0;
      p1_a_sign__1 <= 1'h0;
      p1_or_600 <= 1'h0;
      p2_eq_597 <= 1'h0;
      p2_sel_625 <= 32'h0000_0000;
      p2_not_626 <= 1'h0;
      p2_a_sign__1 <= 1'h0;
      p2_or_600 <= 1'h0;
      p3_a_sign__1 <= 1'h0;
      p3_result <= 32'h0000_0000;
      p0_valid <= 1'h0;
      p1_valid <= 1'h0;
      p2_valid <= 1'h0;
      p3_valid <= 1'h0;
      __xls_float_ips__outs_reg <= 32'h0000_0000;
      __xls_float_ips__outs_valid_reg <= 1'h0;
    end else begin
      p0_a_bexp__2 <= p0_data_enable ? a_bexp__2 : p0_a_bexp__2;
      p0_a_fraction__2 <= p0_data_enable ? a_fraction__2 : p0_a_fraction__2;
      p0_a_sign__1 <= p0_data_enable ? a_sign__1 : p0_a_sign__1;
      p1_a_fraction__2 <= p1_data_enable ? p0_a_fraction__2 : p1_a_fraction__2;
      p1_add_583 <= p1_data_enable ? add_583 : p1_add_583;
      p1_or_594 <= p1_data_enable ? or_594 : p1_or_594;
      p1_eq_597 <= p1_data_enable ? eq_597 : p1_eq_597;
      p1_a_sign__1 <= p1_data_enable ? p0_a_sign__1 : p1_a_sign__1;
      p1_or_600 <= p1_data_enable ? or_600 : p1_or_600;
      p2_eq_597 <= p2_data_enable ? p1_eq_597 : p2_eq_597;
      p2_sel_625 <= p2_data_enable ? sel_625 : p2_sel_625;
      p2_not_626 <= p2_data_enable ? not_626 : p2_not_626;
      p2_a_sign__1 <= p2_data_enable ? p1_a_sign__1 : p2_a_sign__1;
      p2_or_600 <= p2_data_enable ? p1_or_600 : p2_or_600;
      p3_a_sign__1 <= p3_data_enable ? p2_a_sign__1 : p3_a_sign__1;
      p3_result <= p3_data_enable ? result : p3_result;
      p0_valid <= p0_enable ? xls_float_ips__ins_vld : p0_valid;
      p1_valid <= p1_enable ? p0_valid : p1_valid;
      p2_valid <= p2_enable ? p1_valid : p2_valid;
      p3_valid <= p3_enable ? p2_valid : p3_valid;
      __xls_float_ips__outs_reg <= xls_float_ips__outs_load_en ? result__2 : __xls_float_ips__outs_reg;
      __xls_float_ips__outs_valid_reg <= xls_float_ips__outs_valid_load_en ? p3_valid : __xls_float_ips__outs_valid_reg;
    end
  end
  assign xls_float_ips__outs = __xls_float_ips__outs_reg;
  assign xls_float_ips__outs_vld = __xls_float_ips__outs_valid_reg;
  assign xls_float_ips__ins_rdy = p0_data_enable;
endmodule
module __xls_float_ips__mulf32_0_next(
  input wire clk,
  input wire rst,
  input wire [31:0] xls_float_ips__lhs,
  input wire xls_float_ips__lhs_vld,
  input wire [31:0] xls_float_ips__rhs,
  input wire xls_float_ips__rhs_vld,
  input wire xls_float_ips__result_rdy,
  output wire [31:0] xls_float_ips__result,
  output wire xls_float_ips__result_vld,
  output wire xls_float_ips__lhs_rdy,
  output wire xls_float_ips__rhs_rdy
);
  // lint_off MULTIPLY
  function automatic [47:0] umul48b_24b_x_24b (input reg [23:0] lhs, input reg [23:0] rhs);
    begin
      umul48b_24b_x_24b = lhs * rhs;
    end
  endfunction
  // lint_on MULTIPLY
  wire [31:0] __xls_float_ips__result_reg_init = {1'h0, 8'h00, 23'h00_0000};
  reg [47:0] p0_fraction;
  reg p0_bit_slice_907;
  reg p0_bit_slice_908;
  reg [9:0] p0_exp__1;
  reg p0_has_inf_arg;
  reg p0_is_result_nan;
  reg p0_result_sign;
  reg [9:0] p1_exp__2;
  reg [22:0] p1_fraction__5;
  reg p1_greater_than_half_way;
  reg p1_nor_978;
  reg p1_has_inf_arg;
  reg p1_is_result_nan;
  reg p1_result_sign__1;
  reg p2_is_subnormal;
  reg [8:0] p2_result_exp__1;
  reg p2_has_inf_arg;
  reg p2_is_result_nan;
  reg [22:0] p2_result_fraction;
  reg p2_result_sign__1;
  reg p0_valid;
  reg p1_valid;
  reg p2_valid;
  reg [31:0] __xls_float_ips__result_reg;
  reg __xls_float_ips__result_valid_reg;
  wire xls_float_ips__result_valid_inv;
  wire [23:0] fraction__6;
  wire [47:0] fraction__1;
  wire [47:0] sticky;
  wire xls_float_ips__result_valid_load_en;
  wire do_round_up;
  wire [23:0] add_1001;
  wire [47:0] fraction__2;
  wire xls_float_ips__result_load_en;
  wire [23:0] fraction__7;
  wire [9:0] exp__2;
  wire p3_stage_done;
  wire p3_not_valid;
  wire [7:0] a_bexp__3;
  wire [7:0] b_bexp__8;
  wire and_reduce_1030;
  wire [9:0] add_1005;
  wire p2_enable;
  wire eq_883;
  wire eq_884;
  wire [7:0] high_exp;
  wire [22:0] a_fraction__3;
  wire [7:0] high_exp__1;
  wire [22:0] b_fraction__6;
  wire [9:0] exp__3;
  wire [47:0] fraction__3;
  wire [47:0] sticky__1;
  wire p2_data_enable;
  wire p2_not_valid;
  wire eq_916;
  wire eq_917;
  wire eq_918;
  wire eq_919;
  wire is_subnormal;
  wire [47:0] fraction__4;
  wire p1_enable;
  wire [8:0] add_902;
  wire p1_data_enable;
  wire p1_not_valid;
  wire [23:0] a_fraction__1;
  wire [23:0] b_fraction__1;
  wire has_0_arg;
  wire has_inf_arg;
  wire [7:0] high_exp__2;
  wire [22:0] result_fraction__3;
  wire [22:0] nan_fraction;
  wire [8:0] result_exp;
  wire ne_973;
  wire p0_enable;
  wire p0_all_active_inputs_valid;
  wire [47:0] fraction;
  wire [9:0] exp;
  wire a_sign__1;
  wire b_sign__1;
  wire [7:0] result_exp__4;
  wire [22:0] result_fraction__4;
  wire [8:0] result_exp__1;
  wire [22:0] result_fraction;
  wire [22:0] fraction__5;
  wire greater_than_half_way;
  wire nor_978;
  wire result_sign__1;
  wire p0_data_enable;
  wire bit_slice_907;
  wire bit_slice_908;
  wire [9:0] exp__1;
  wire is_result_nan;
  wire result_sign;
  wire [31:0] __xls_float_ips__result_buf;
  assign xls_float_ips__result_valid_inv = ~__xls_float_ips__result_valid_reg;
  assign fraction__6 = {1'h0, p1_fraction__5};
  assign fraction__1 = p0_fraction >> p0_bit_slice_907;
  assign sticky = {47'h0000_0000_0000, p0_bit_slice_908};
  assign xls_float_ips__result_valid_load_en = xls_float_ips__result_rdy | xls_float_ips__result_valid_inv;
  assign do_round_up = p1_greater_than_half_way | p1_nor_978;
  assign add_1001 = fraction__6 + 24'h00_0001;
  assign fraction__2 = fraction__1 | sticky;
  assign xls_float_ips__result_load_en = p2_valid & xls_float_ips__result_valid_load_en;
  assign fraction__7 = do_round_up ? add_1001 : fraction__6;
  assign exp__2 = p0_exp__1 + {9'h000, p0_bit_slice_907};
  assign p3_stage_done = p2_valid & xls_float_ips__result_load_en;
  assign p3_not_valid = ~p2_valid;
  assign a_bexp__3 = xls_float_ips__lhs[30:23];
  assign b_bexp__8 = xls_float_ips__rhs[30:23];
  assign and_reduce_1030 = &p2_result_exp__1[7:0];
  assign add_1005 = p1_exp__2 + 10'h001;
  assign p2_enable = p3_stage_done | p3_not_valid;
  assign eq_883 = a_bexp__3 == 8'h00;
  assign eq_884 = b_bexp__8 == 8'h00;
  assign high_exp = 8'hff;
  assign a_fraction__3 = xls_float_ips__lhs[22:0];
  assign high_exp__1 = 8'hff;
  assign b_fraction__6 = xls_float_ips__rhs[22:0];
  assign exp__3 = fraction__7[23] ? add_1005 : p1_exp__2;
  assign fraction__3 = $signed(exp__2) <= $signed(10'h000) ? {1'h0, fraction__2[47:1]} : fraction__2;
  assign sticky__1 = {47'h0000_0000_0000, fraction__2[0]};
  assign p2_data_enable = p2_enable & p1_valid;
  assign p2_not_valid = ~p1_valid;
  assign eq_916 = a_bexp__3 == high_exp;
  assign eq_917 = a_fraction__3 == 23'h00_0000;
  assign eq_918 = b_bexp__8 == high_exp__1;
  assign eq_919 = b_fraction__6 == 23'h00_0000;
  assign is_subnormal = $signed(exp__3) <= $signed(10'h000);
  assign fraction__4 = fraction__3 | sticky__1;
  assign p1_enable = p2_data_enable | p2_not_valid;
  assign add_902 = {1'h0, a_bexp__3} + {1'h0, b_bexp__8};
  assign p1_data_enable = p1_enable & p0_valid;
  assign p1_not_valid = ~p0_valid;
  assign a_fraction__1 = {1'h1, a_fraction__3} & {24{~eq_883}};
  assign b_fraction__1 = {1'h1, b_fraction__6} & {24{~eq_884}};
  assign has_0_arg = eq_883 | eq_884;
  assign has_inf_arg = eq_916 & eq_917 | eq_918 & eq_919;
  assign high_exp__2 = 8'hff;
  assign result_fraction__3 = p2_result_fraction & {23{~(p2_has_inf_arg | p2_result_exp__1[8] | and_reduce_1030 | p2_is_subnormal)}};
  assign nan_fraction = 23'h40_0000;
  assign result_exp = exp__3[8:0];
  assign ne_973 = fraction__4[21:0] != 22'h00_0000;
  assign p0_enable = p1_data_enable | p1_not_valid;
  assign p0_all_active_inputs_valid = xls_float_ips__lhs_vld & xls_float_ips__rhs_vld;
  assign fraction = umul48b_24b_x_24b(a_fraction__1, b_fraction__1);
  assign exp = {1'h0, add_902} + 10'h381;
  assign a_sign__1 = xls_float_ips__lhs[31:31];
  assign b_sign__1 = xls_float_ips__rhs[31:31];
  assign result_exp__4 = p2_is_result_nan | p2_has_inf_arg | p2_result_exp__1[8] | and_reduce_1030 ? high_exp__2 : p2_result_exp__1[7:0];
  assign result_fraction__4 = p2_is_result_nan ? nan_fraction : result_fraction__3;
  assign result_exp__1 = result_exp & {9{~is_subnormal}};
  assign result_fraction = fraction__7[22:0];
  assign fraction__5 = fraction__4[45:23];
  assign greater_than_half_way = fraction__4[22] & ne_973;
  assign nor_978 = ~(~fraction__4[22] | ne_973 | ~fraction__4[23]);
  assign result_sign__1 = ~p0_is_result_nan & p0_result_sign;
  assign p0_data_enable = p0_enable & p0_all_active_inputs_valid;
  assign bit_slice_907 = fraction[47];
  assign bit_slice_908 = fraction[0];
  assign exp__1 = exp & {10{~(eq_883 | eq_884)}};
  assign is_result_nan = ~(~eq_916 | eq_917) | ~(~eq_918 | eq_919) | has_0_arg & has_inf_arg;
  assign result_sign = a_sign__1 ^ b_sign__1;
  assign __xls_float_ips__result_buf = {p2_result_sign__1, result_exp__4, result_fraction__4};
  always @ (posedge clk) begin
    if (rst) begin
      p0_fraction <= 48'h0000_0000_0000;
      p0_bit_slice_907 <= 1'h0;
      p0_bit_slice_908 <= 1'h0;
      p0_exp__1 <= 10'h000;
      p0_has_inf_arg <= 1'h0;
      p0_is_result_nan <= 1'h0;
      p0_result_sign <= 1'h0;
      p1_exp__2 <= 10'h000;
      p1_fraction__5 <= 23'h00_0000;
      p1_greater_than_half_way <= 1'h0;
      p1_nor_978 <= 1'h0;
      p1_has_inf_arg <= 1'h0;
      p1_is_result_nan <= 1'h0;
      p1_result_sign__1 <= 1'h0;
      p2_is_subnormal <= 1'h0;
      p2_result_exp__1 <= 9'h000;
      p2_has_inf_arg <= 1'h0;
      p2_is_result_nan <= 1'h0;
      p2_result_fraction <= 23'h00_0000;
      p2_result_sign__1 <= 1'h0;
      p0_valid <= 1'h0;
      p1_valid <= 1'h0;
      p2_valid <= 1'h0;
      __xls_float_ips__result_reg <= __xls_float_ips__result_reg_init;
      __xls_float_ips__result_valid_reg <= 1'h0;
    end else begin
      p0_fraction <= p0_data_enable ? fraction : p0_fraction;
      p0_bit_slice_907 <= p0_data_enable ? bit_slice_907 : p0_bit_slice_907;
      p0_bit_slice_908 <= p0_data_enable ? bit_slice_908 : p0_bit_slice_908;
      p0_exp__1 <= p0_data_enable ? exp__1 : p0_exp__1;
      p0_has_inf_arg <= p0_data_enable ? has_inf_arg : p0_has_inf_arg;
      p0_is_result_nan <= p0_data_enable ? is_result_nan : p0_is_result_nan;
      p0_result_sign <= p0_data_enable ? result_sign : p0_result_sign;
      p1_exp__2 <= p1_data_enable ? exp__2 : p1_exp__2;
      p1_fraction__5 <= p1_data_enable ? fraction__5 : p1_fraction__5;
      p1_greater_than_half_way <= p1_data_enable ? greater_than_half_way : p1_greater_than_half_way;
      p1_nor_978 <= p1_data_enable ? nor_978 : p1_nor_978;
      p1_has_inf_arg <= p1_data_enable ? p0_has_inf_arg : p1_has_inf_arg;
      p1_is_result_nan <= p1_data_enable ? p0_is_result_nan : p1_is_result_nan;
      p1_result_sign__1 <= p1_data_enable ? result_sign__1 : p1_result_sign__1;
      p2_is_subnormal <= p2_data_enable ? is_subnormal : p2_is_subnormal;
      p2_result_exp__1 <= p2_data_enable ? result_exp__1 : p2_result_exp__1;
      p2_has_inf_arg <= p2_data_enable ? p1_has_inf_arg : p2_has_inf_arg;
      p2_is_result_nan <= p2_data_enable ? p1_is_result_nan : p2_is_result_nan;
      p2_result_fraction <= p2_data_enable ? result_fraction : p2_result_fraction;
      p2_result_sign__1 <= p2_data_enable ? p1_result_sign__1 : p2_result_sign__1;
      p0_valid <= p0_enable ? p0_all_active_inputs_valid : p0_valid;
      p1_valid <= p1_enable ? p0_valid : p1_valid;
      p2_valid <= p2_enable ? p1_valid : p2_valid;
      __xls_float_ips__result_reg <= xls_float_ips__result_load_en ? __xls_float_ips__result_buf : __xls_float_ips__result_reg;
      __xls_float_ips__result_valid_reg <= xls_float_ips__result_valid_load_en ? p2_valid : __xls_float_ips__result_valid_reg;
    end
  end
  assign xls_float_ips__result = __xls_float_ips__result_reg;
  assign xls_float_ips__result_vld = __xls_float_ips__result_valid_reg;
  assign xls_float_ips__lhs_rdy = p0_data_enable;
  assign xls_float_ips__rhs_rdy = p0_data_enable;
endmodule
module __xls_float_ips__sitofp_0_next(
  input wire clk,
  input wire rst,
  input wire [31:0] xls_float_ips__ins,
  input wire xls_float_ips__ins_vld,
  input wire xls_float_ips__outs_rdy,
  output wire [31:0] xls_float_ips__outs,
  output wire xls_float_ips__outs_vld,
  output wire xls_float_ips__ins_rdy
);
  wire [31:0] __xls_float_ips__outs_reg_init = {1'h0, 8'h00, 23'h00_0000};
  reg p0_sign;
  reg [30:0] p0_fraction;
  reg [30:0] p0_reverse_395;
  reg p0_is_neg_int_max;
  reg p1_sign;
  reg [4:0] p1_encode_411;
  reg [6:0] p1_bit_slice_418;
  reg [25:0] p1_bit_slice_419;
  reg p1_is_neg_int_max;
  reg p2_sign;
  reg [23:0] p2_concat_448;
  reg p2_do_round_up;
  reg [23:0] p2_add_452;
  reg [7:0] p2_bexp;
  reg p2_is_neg_int_max;
  reg p3_sign;
  reg [7:0] p3_bexp__1;
  reg [22:0] p3_fraction__4;
  reg p3_is_neg_int_max;
  reg p3_nor_481;
  reg p3_or_482;
  reg p0_valid;
  reg p1_valid;
  reg p2_valid;
  reg p3_valid;
  reg [31:0] __xls_float_ips__outs_reg;
  reg __xls_float_ips__outs_valid_reg;
  wire xls_float_ips__outs_valid_inv;
  wire xls_float_ips__outs_valid_load_en;
  wire xls_float_ips__outs_load_en;
  wire p4_stage_done;
  wire p4_not_valid;
  wire p3_enable;
  wire p3_data_enable;
  wire p3_not_valid;
  wire [23:0] fraction__3_squeezed_portion_3_width_24;
  wire [31:0] one_hot_409;
  wire p2_enable;
  wire [7:0] add_473;
  wire [4:0] encode_411;
  wire p2_data_enable;
  wire p2_not_valid;
  wire [7:0] bexp__1;
  wire [25:0] fraction__2;
  wire p1_enable;
  wire [22:0] fraction__4;
  wire [2:0] normal_chunk;
  wire [1:0] half_way_chunk;
  wire [6:0] sub_450;
  wire [5:0] add_416;
  wire p1_data_enable;
  wire p1_not_valid;
  wire sign;
  wire and_reduce_479;
  wire ne_480;
  wire [23:0] concat_448;
  wire [7:0] exp;
  wire [32:0] fraction__1;
  wire p0_enable;
  wire [30:0] fraction;
  wire nor_481;
  wire or_482;
  wire do_round_up;
  wire [23:0] add_452;
  wire [7:0] bexp;
  wire [6:0] bit_slice_418;
  wire [25:0] bit_slice_419;
  wire p0_data_enable;
  wire [30:0] reverse_395;
  wire is_neg_int_max;
  wire [31:0] result__2;
  assign xls_float_ips__outs_valid_inv = ~__xls_float_ips__outs_valid_reg;
  assign xls_float_ips__outs_valid_load_en = xls_float_ips__outs_rdy | xls_float_ips__outs_valid_inv;
  assign xls_float_ips__outs_load_en = p3_valid & xls_float_ips__outs_valid_load_en;
  assign p4_stage_done = p3_valid & xls_float_ips__outs_load_en;
  assign p4_not_valid = ~p3_valid;
  assign p3_enable = p4_stage_done | p4_not_valid;
  assign p3_data_enable = p3_enable & p2_valid;
  assign p3_not_valid = ~p2_valid;
  assign fraction__3_squeezed_portion_3_width_24 = p2_do_round_up ? p2_add_452 : p2_concat_448;
  assign one_hot_409 = {p0_reverse_395[30:0] == 31'h0000_0000, p0_reverse_395[30] && p0_reverse_395[29:0] == 30'h0000_0000, p0_reverse_395[29] && p0_reverse_395[28:0] == 29'h0000_0000, p0_reverse_395[28] && p0_reverse_395[27:0] == 28'h000_0000, p0_reverse_395[27] && p0_reverse_395[26:0] == 27'h000_0000, p0_reverse_395[26] && p0_reverse_395[25:0] == 26'h000_0000, p0_reverse_395[25] && p0_reverse_395[24:0] == 25'h000_0000, p0_reverse_395[24] && p0_reverse_395[23:0] == 24'h00_0000, p0_reverse_395[23] && p0_reverse_395[22:0] == 23'h00_0000, p0_reverse_395[22] && p0_reverse_395[21:0] == 22'h00_0000, p0_reverse_395[21] && p0_reverse_395[20:0] == 21'h00_0000, p0_reverse_395[20] && p0_reverse_395[19:0] == 20'h0_0000, p0_reverse_395[19] && p0_reverse_395[18:0] == 19'h0_0000, p0_reverse_395[18] && p0_reverse_395[17:0] == 18'h0_0000, p0_reverse_395[17] && p0_reverse_395[16:0] == 17'h0_0000, p0_reverse_395[16] && p0_reverse_395[15:0] == 16'h0000, p0_reverse_395[15] && p0_reverse_395[14:0] == 15'h0000, p0_reverse_395[14] && p0_reverse_395[13:0] == 14'h0000, p0_reverse_395[13] && p0_reverse_395[12:0] == 13'h0000, p0_reverse_395[12] && p0_reverse_395[11:0] == 12'h000, p0_reverse_395[11] && p0_reverse_395[10:0] == 11'h000, p0_reverse_395[10] && p0_reverse_395[9:0] == 10'h000, p0_reverse_395[9] && p0_reverse_395[8:0] == 9'h000, p0_reverse_395[8] && p0_reverse_395[7:0] == 8'h00, p0_reverse_395[7] && p0_reverse_395[6:0] == 7'h00, p0_reverse_395[6] && p0_reverse_395[5:0] == 6'h00, p0_reverse_395[5] && p0_reverse_395[4:0] == 5'h00, p0_reverse_395[4] && p0_reverse_395[3:0] == 4'h0, p0_reverse_395[3] && p0_reverse_395[2:0] == 3'h0, p0_reverse_395[2] && p0_reverse_395[1:0] == 2'h0, p0_reverse_395[1] && !p0_reverse_395[0], p0_reverse_395[0]};
  assign p2_enable = p3_data_enable | p3_not_valid;
  assign add_473 = p2_bexp + 8'h01;
  assign encode_411 = {one_hot_409[16] | one_hot_409[17] | one_hot_409[18] | one_hot_409[19] | one_hot_409[20] | one_hot_409[21] | one_hot_409[22] | one_hot_409[23] | one_hot_409[24] | one_hot_409[25] | one_hot_409[26] | one_hot_409[27] | one_hot_409[28] | one_hot_409[29] | one_hot_409[30] | one_hot_409[31], one_hot_409[8] | one_hot_409[9] | one_hot_409[10] | one_hot_409[11] | one_hot_409[12] | one_hot_409[13] | one_hot_409[14] | one_hot_409[15] | one_hot_409[24] | one_hot_409[25] | one_hot_409[26] | one_hot_409[27] | one_hot_409[28] | one_hot_409[29] | one_hot_409[30] | one_hot_409[31], one_hot_409[4] | one_hot_409[5] | one_hot_409[6] | one_hot_409[7] | one_hot_409[12] | one_hot_409[13] | one_hot_409[14] | one_hot_409[15] | one_hot_409[20] | one_hot_409[21] | one_hot_409[22] | one_hot_409[23] | one_hot_409[28] | one_hot_409[29] | one_hot_409[30] | one_hot_409[31], one_hot_409[2] | one_hot_409[3] | one_hot_409[6] | one_hot_409[7] | one_hot_409[10] | one_hot_409[11] | one_hot_409[14] | one_hot_409[15] | one_hot_409[18] | one_hot_409[19] | one_hot_409[22] | one_hot_409[23] | one_hot_409[26] | one_hot_409[27] | one_hot_409[30] | one_hot_409[31], one_hot_409[1] | one_hot_409[3] | one_hot_409[5] | one_hot_409[7] | one_hot_409[9] | one_hot_409[11] | one_hot_409[13] | one_hot_409[15] | one_hot_409[17] | one_hot_409[19] | one_hot_409[21] | one_hot_409[23] | one_hot_409[25] | one_hot_409[27] | one_hot_409[29] | one_hot_409[31]};
  assign p2_data_enable = p2_enable & p1_valid;
  assign p2_not_valid = ~p1_valid;
  assign bexp__1 = fraction__3_squeezed_portion_3_width_24[23] ? add_473 : p2_bexp;
  assign fraction__2 = p1_bit_slice_419 | {25'h000_0000, p1_bit_slice_418 != 7'h00};
  assign p1_enable = p2_data_enable | p2_not_valid;
  assign fraction__4 = fraction__3_squeezed_portion_3_width_24[22:0];
  assign normal_chunk = fraction__2[2:0];
  assign half_way_chunk = fraction__2[3:2];
  assign sub_450 = 7'h1e - {2'h0, p1_encode_411};
  assign add_416 = {1'h0, encode_411} + 6'h03;
  assign p1_data_enable = p1_enable & p0_valid;
  assign p1_not_valid = ~p0_valid;
  assign sign = xls_float_ips__ins[31];
  assign and_reduce_479 = &bexp__1[6:0];
  assign ne_480 = fraction__4 != 23'h00_0000;
  assign concat_448 = {1'h0, fraction__2[25:3]};
  assign exp = {{1{sub_450[6]}}, sub_450};
  assign fraction__1 = add_416 >= 6'h21 ? 33'h0_0000_0000 : {2'h0, p0_fraction} << add_416;
  assign p0_enable = p1_data_enable | p1_not_valid;
  assign fraction = sign ? -xls_float_ips__ins[30:0] : xls_float_ips__ins[30:0];
  assign nor_481 = ~(bexp__1[7] | and_reduce_479 | ne_480);
  assign or_482 = bexp__1[7] | and_reduce_479 | ne_480;
  assign do_round_up = normal_chunk > 3'h4 | half_way_chunk == 2'h3;
  assign add_452 = concat_448 + 24'h00_0001;
  assign bexp = exp + 8'h7f;
  assign bit_slice_418 = fraction__1[6:0];
  assign bit_slice_419 = fraction__1[32:7];
  assign p0_data_enable = p0_enable & xls_float_ips__ins_vld;
  assign reverse_395 = {fraction[0], fraction[1], fraction[2], fraction[3], fraction[4], fraction[5], fraction[6], fraction[7], fraction[8], fraction[9], fraction[10], fraction[11], fraction[12], fraction[13], fraction[14], fraction[15], fraction[16], fraction[17], fraction[18], fraction[19], fraction[20], fraction[21], fraction[22], fraction[23], fraction[24], fraction[25], fraction[26], fraction[27], fraction[28], fraction[29], fraction[30]};
  assign is_neg_int_max = xls_float_ips__ins == 32'h8000_0000;
  assign result__2 = {p3_is_neg_int_max | ~p3_is_neg_int_max & p3_or_482 & p3_sign, p3_is_neg_int_max ? 8'h9e : p3_bexp__1 & {8{p3_or_482}}, p3_fraction__4 & {23{~(p3_is_neg_int_max | p3_nor_481)}}};
  always @ (posedge clk) begin
    if (rst) begin
      p0_sign <= 1'h0;
      p0_fraction <= 31'h0000_0000;
      p0_reverse_395 <= 31'h0000_0000;
      p0_is_neg_int_max <= 1'h0;
      p1_sign <= 1'h0;
      p1_encode_411 <= 5'h00;
      p1_bit_slice_418 <= 7'h00;
      p1_bit_slice_419 <= 26'h000_0000;
      p1_is_neg_int_max <= 1'h0;
      p2_sign <= 1'h0;
      p2_concat_448 <= 24'h00_0000;
      p2_do_round_up <= 1'h0;
      p2_add_452 <= 24'h00_0000;
      p2_bexp <= 8'h00;
      p2_is_neg_int_max <= 1'h0;
      p3_sign <= 1'h0;
      p3_bexp__1 <= 8'h00;
      p3_fraction__4 <= 23'h00_0000;
      p3_is_neg_int_max <= 1'h0;
      p3_nor_481 <= 1'h0;
      p3_or_482 <= 1'h0;
      p0_valid <= 1'h0;
      p1_valid <= 1'h0;
      p2_valid <= 1'h0;
      p3_valid <= 1'h0;
      __xls_float_ips__outs_reg <= __xls_float_ips__outs_reg_init;
      __xls_float_ips__outs_valid_reg <= 1'h0;
    end else begin
      p0_sign <= p0_data_enable ? sign : p0_sign;
      p0_fraction <= p0_data_enable ? fraction : p0_fraction;
      p0_reverse_395 <= p0_data_enable ? reverse_395 : p0_reverse_395;
      p0_is_neg_int_max <= p0_data_enable ? is_neg_int_max : p0_is_neg_int_max;
      p1_sign <= p1_data_enable ? p0_sign : p1_sign;
      p1_encode_411 <= p1_data_enable ? encode_411 : p1_encode_411;
      p1_bit_slice_418 <= p1_data_enable ? bit_slice_418 : p1_bit_slice_418;
      p1_bit_slice_419 <= p1_data_enable ? bit_slice_419 : p1_bit_slice_419;
      p1_is_neg_int_max <= p1_data_enable ? p0_is_neg_int_max : p1_is_neg_int_max;
      p2_sign <= p2_data_enable ? p1_sign : p2_sign;
      p2_concat_448 <= p2_data_enable ? concat_448 : p2_concat_448;
      p2_do_round_up <= p2_data_enable ? do_round_up : p2_do_round_up;
      p2_add_452 <= p2_data_enable ? add_452 : p2_add_452;
      p2_bexp <= p2_data_enable ? bexp : p2_bexp;
      p2_is_neg_int_max <= p2_data_enable ? p1_is_neg_int_max : p2_is_neg_int_max;
      p3_sign <= p3_data_enable ? p2_sign : p3_sign;
      p3_bexp__1 <= p3_data_enable ? bexp__1 : p3_bexp__1;
      p3_fraction__4 <= p3_data_enable ? fraction__4 : p3_fraction__4;
      p3_is_neg_int_max <= p3_data_enable ? p2_is_neg_int_max : p3_is_neg_int_max;
      p3_nor_481 <= p3_data_enable ? nor_481 : p3_nor_481;
      p3_or_482 <= p3_data_enable ? or_482 : p3_or_482;
      p0_valid <= p0_enable ? xls_float_ips__ins_vld : p0_valid;
      p1_valid <= p1_enable ? p0_valid : p1_valid;
      p2_valid <= p2_enable ? p1_valid : p2_valid;
      p3_valid <= p3_enable ? p2_valid : p3_valid;
      __xls_float_ips__outs_reg <= xls_float_ips__outs_load_en ? result__2 : __xls_float_ips__outs_reg;
      __xls_float_ips__outs_valid_reg <= xls_float_ips__outs_valid_load_en ? p3_valid : __xls_float_ips__outs_valid_reg;
    end
  end
  assign xls_float_ips__outs = __xls_float_ips__outs_reg;
  assign xls_float_ips__outs_vld = __xls_float_ips__outs_valid_reg;
  assign xls_float_ips__ins_rdy = p0_data_enable;
endmodule
module __xls_float_ips__subf32_0_next(
  input wire clk,
  input wire rst,
  input wire [31:0] xls_float_ips__rhs,
  input wire xls_float_ips__rhs_vld,
  input wire [31:0] xls_float_ips__lhs,
  input wire xls_float_ips__lhs_vld,
  input wire xls_float_ips__result_rdy,
  output wire [31:0] xls_float_ips__result,
  output wire xls_float_ips__result_vld,
  output wire xls_float_ips__rhs_rdy,
  output wire xls_float_ips__lhs_rdy
);
  function automatic [3:0] priority_sel_4b_2way (input reg [1:0] sel, input reg [3:0] case0, input reg [3:0] case1, input reg [3:0] default_value);
    begin
      casez (sel)
        2'b?1: begin
          priority_sel_4b_2way = case0;
        end
        2'b10: begin
          priority_sel_4b_2way = case1;
        end
        2'b00: begin
          priority_sel_4b_2way = default_value;
        end
        default: begin
          // Propagate X
          priority_sel_4b_2way = 4'dx;
        end
      endcase
    end
  endfunction
  function automatic [1:0] priority_sel_2b_2way (input reg [1:0] sel, input reg [1:0] case0, input reg [1:0] case1, input reg [1:0] default_value);
    begin
      casez (sel)
        2'b?1: begin
          priority_sel_2b_2way = case0;
        end
        2'b10: begin
          priority_sel_2b_2way = case1;
        end
        2'b00: begin
          priority_sel_2b_2way = default_value;
        end
        default: begin
          // Propagate X
          priority_sel_2b_2way = 2'dx;
        end
      endcase
    end
  endfunction
  function automatic priority_sel_1b_4way (input reg [3:0] sel, input reg case0, input reg case1, input reg case2, input reg case3, input reg default_value);
    begin
      casez (sel)
        4'b???1: begin
          priority_sel_1b_4way = case0;
        end
        4'b??10: begin
          priority_sel_1b_4way = case1;
        end
        4'b?100: begin
          priority_sel_1b_4way = case2;
        end
        4'b1000: begin
          priority_sel_1b_4way = case3;
        end
        4'b0000: begin
          priority_sel_1b_4way = default_value;
        end
        default: begin
          // Propagate X
          priority_sel_1b_4way = 1'dx;
        end
      endcase
    end
  endfunction
  function automatic priority_sel_1b_3way (input reg [2:0] sel, input reg case0, input reg case1, input reg case2, input reg default_value);
    begin
      casez (sel)
        3'b??1: begin
          priority_sel_1b_3way = case0;
        end
        3'b?10: begin
          priority_sel_1b_3way = case1;
        end
        3'b100: begin
          priority_sel_1b_3way = case2;
        end
        3'b000: begin
          priority_sel_1b_3way = default_value;
        end
        default: begin
          // Propagate X
          priority_sel_1b_3way = 1'dx;
        end
      endcase
    end
  endfunction
  function automatic [2:0] priority_sel_3b_2way (input reg [1:0] sel, input reg [2:0] case0, input reg [2:0] case1, input reg [2:0] default_value);
    begin
      casez (sel)
        2'b?1: begin
          priority_sel_3b_2way = case0;
        end
        2'b10: begin
          priority_sel_3b_2way = case1;
        end
        2'b00: begin
          priority_sel_3b_2way = default_value;
        end
        default: begin
          // Propagate X
          priority_sel_3b_2way = 3'dx;
        end
      endcase
    end
  endfunction
  function automatic [1:0] priority_sel_2b_4way (input reg [3:0] sel, input reg [1:0] case0, input reg [1:0] case1, input reg [1:0] case2, input reg [1:0] case3, input reg [1:0] default_value);
    begin
      casez (sel)
        4'b???1: begin
          priority_sel_2b_4way = case0;
        end
        4'b??10: begin
          priority_sel_2b_4way = case1;
        end
        4'b?100: begin
          priority_sel_2b_4way = case2;
        end
        4'b1000: begin
          priority_sel_2b_4way = case3;
        end
        4'b0000: begin
          priority_sel_2b_4way = default_value;
        end
        default: begin
          // Propagate X
          priority_sel_2b_4way = 2'dx;
        end
      endcase
    end
  endfunction
  function automatic priority_sel_1b_2way (input reg [1:0] sel, input reg case0, input reg case1, input reg default_value);
    begin
      casez (sel)
        2'b?1: begin
          priority_sel_1b_2way = case0;
        end
        2'b10: begin
          priority_sel_1b_2way = case1;
        end
        2'b00: begin
          priority_sel_1b_2way = default_value;
        end
        default: begin
          // Propagate X
          priority_sel_1b_2way = 1'dx;
        end
      endcase
    end
  endfunction
  wire [31:0] __xls_float_ips__result_reg_init = {1'h0, 8'h00, 23'h00_0000};
  reg [7:0] p0_b_bexp__6;
  reg [7:0] p0_a_bexp__2;
  reg p0_bit_slice_107413;
  reg [22:0] p0_b_fraction__6;
  reg [22:0] p0_tuple_index_107415;
  reg [7:0] p0_bit_slice_107416;
  reg p0_not_107418;
  reg p0_tuple_index_107419;
  reg [7:0] p1_a_bexp__4;
  reg p1_b_sign__3;
  reg p1_xor_107473;
  reg [24:0] p1_wide_x_squeezed;
  reg [24:0] p1_bit_slice_107475;
  reg [27:0] p1_shrl_107476;
  reg p1_sticky;
  reg p1_is_operand_inf;
  reg p1_and_107506;
  reg p1_is_result_nan;
  reg p1_not_107508;
  reg [7:0] p2_a_bexp__4;
  reg [27:0] p2_abs_fraction__1;
  reg p2_not_107554;
  reg p2_is_operand_inf;
  reg p2_is_result_nan;
  reg p2_result_sign;
  reg p2_not_107508;
  reg [7:0] p3_a_bexp__4;
  reg [27:0] p3_abs_fraction__1;
  reg p3_carry_bit;
  reg p3_and_107695;
  reg p3_and_107697;
  reg p3_nor_107703;
  reg p3_nor_107730;
  reg p3_leading_zeroes__4_to_5;
  reg [2:0] p3_priority_sel_107732;
  reg [1:0] p3_priority_sel_107733;
  reg [2:0] p3_priority_sel_107734;
  reg p3_or_107735;
  reg p3_not_107554;
  reg p3_is_operand_inf;
  reg p3_is_result_nan;
  reg p3_result_sign__2;
  reg [7:0] p4_a_bexp__4;
  reg p4_leading_zeroes__4_to_5;
  reg [3:0] p4_leading_zeroes__0_to_4;
  reg [2:0] p4_normal_chunk;
  reg [1:0] p4_half_way_chunk;
  reg [23:0] p4_bit_slice_107789;
  reg p4_not_107554;
  reg p4_is_operand_inf;
  reg p4_is_result_nan;
  reg p4_result_sign__2;
  reg p5_leading_zeroes__4_to_5;
  reg [3:0] p5_leading_zeroes__0_to_4;
  reg [9:0] p5_concat_107829;
  reg p5_not_107554;
  reg p5_is_operand_inf;
  reg p5_is_result_nan;
  reg [22:0] p5_result_fraction;
  reg p5_result_sign__2;
  reg [8:0] p6_wide_exponent__2;
  reg p6_is_operand_inf;
  reg p6_is_result_nan;
  reg [22:0] p6_result_fraction;
  reg p6_result_sign__2;
  reg p7_is_result_nan;
  reg [22:0] p7_result_fraction__3;
  reg p7_result_sign__2;
  reg [7:0] p7_result_exponent__2;
  reg p0_valid;
  reg p1_valid;
  reg p2_valid;
  reg p3_valid;
  reg p4_valid;
  reg p5_valid;
  reg p6_valid;
  reg p7_valid;
  reg [31:0] __xls_float_ips__result_reg;
  reg __xls_float_ips__result_valid_reg;
  wire xls_float_ips__result_valid_inv;
  wire xls_float_ips__result_valid_load_en;
  wire xls_float_ips__result_load_en;
  wire p8_stage_done;
  wire p8_not_valid;
  wire p7_enable;
  wire p7_data_enable;
  wire p7_not_valid;
  wire p6_enable;
  wire p6_data_enable;
  wire p6_not_valid;
  wire p5_enable;
  wire p5_data_enable;
  wire p5_not_valid;
  wire p4_enable;
  wire p4_data_enable;
  wire p4_not_valid;
  wire [2:0] fraction_shift__3;
  wire p3_enable;
  wire [9:0] add_107856;
  wire [24:0] concat_107817;
  wire carry_bit;
  wire [24:0] addend_x__2_squeezed;
  wire [7:0] a_bexp__4;
  wire [7:0] incremented_sum__1;
  wire [7:0] MAX_EXPONENT;
  wire [22:0] a_fraction__1;
  wire [7:0] b_bexp__7;
  wire [7:0] MAX_EXPONENT__1;
  wire [22:0] b_fraction__7;
  wire p3_data_enable;
  wire p3_not_valid;
  wire [9:0] wide_exponent;
  wire do_round_up;
  wire [24:0] add_107820;
  wire [3:0] leading_zeroes__0_to_4;
  wire nor_107602;
  wire nor_107603;
  wire nor_107605;
  wire nor_107606;
  wire nor_107611;
  wire nor_107612;
  wire nor_107617;
  wire nor_107620;
  wire nor_107621;
  wire nor_107622;
  wire nor_107628;
  wire [7:0] a_bexpbs_difference__2;
  wire eq_107486;
  wire eq_107487;
  wire eq_107488;
  wire eq_107489;
  wire p2_enable;
  wire and_reduce_107883;
  wire [9:0] wide_exponent__1;
  wire [24:0] rounded_fraction_squeezed_portion_3_width_25;
  wire [4:0] leading_zeroes;
  wire nor_107629;
  wire and_107630;
  wire and_107632;
  wire nor_107637;
  wire and_107638;
  wire nor_107641;
  wire and_107645;
  wire nor_107646;
  wire and_107650;
  wire nor_107652;
  wire [25:0] add_107538;
  wire [23:0] fraction_x;
  wire a_sign__1;
  wire b_sign__3;
  wire p2_data_enable;
  wire p2_not_valid;
  wire [7:0] b_bexp__6;
  wire rounding_carry;
  wire [2:0] fraction_shift__2;
  wire [2:0] fraction_shift__4;
  wire [28:0] cancel_fraction;
  wire and_107659;
  wire and_107677;
  wire [23:0] fraction_x__1;
  wire [2:0] addend_x__2_squeezed_const_lsb_bits__1;
  wire [23:0] fraction_y;
  wire [23:0] sign_ext_107458;
  wire [27:0] add_107477;
  wire p1_enable;
  wire [7:0] a_bexp__2;
  wire [27:0] rounded_fraction;
  wire [2:0] fraction_shift__1;
  wire [26:0] cancel_fraction__1;
  wire [26:0] carry_fraction__1;
  wire and_107695;
  wire and_107697;
  wire nor_107703;
  wire and_107704;
  wire [1:0] priority_sel_107711;
  wire [27:0] concat_107543;
  wire fraction_is_zero;
  wire [27:0] wide_x;
  wire [23:0] fraction_y__1;
  wire [2:0] addend_x__2_squeezed_const_lsb_bits;
  wire has_pos_inf;
  wire has_neg_inf;
  wire p1_data_enable;
  wire p1_not_valid;
  wire [22:0] FRACTION_HIGH_BIT;
  wire [22:0] sign_ext_107887;
  wire [7:0] MAX_EXPONENT__2;
  wire [8:0] add_107828;
  wire [27:0] shrl_107834;
  wire [26:0] shifted_fraction;
  wire [2:0] concat_107717;
  wire [2:0] concat_107718;
  wire [2:0] concat_107719;
  wire [1:0] concat_107722;
  wire [2:0] concat_107728;
  wire result_sign__1;
  wire [27:0] neg_107469;
  wire [27:0] wide_y;
  wire p0_enable;
  wire p0_all_active_inputs_valid;
  wire [8:0] sum;
  wire b_sign__2;
  wire [22:0] result_fraction__4;
  wire [22:0] result_fraction__3;
  wire [7:0] result_exponent__2;
  wire [8:0] wide_exponent__2;
  wire [9:0] concat_107829;
  wire [22:0] result_fraction;
  wire [2:0] normal_chunk;
  wire [1:0] half_way_chunk;
  wire [23:0] bit_slice_107789;
  wire nor_107730;
  wire leading_zeroes__4_to_5;
  wire [2:0] priority_sel_107732;
  wire [1:0] priority_sel_107733;
  wire [2:0] priority_sel_107734;
  wire or_107735;
  wire result_sign__2;
  wire [27:0] abs_fraction__1;
  wire not_107554;
  wire result_sign;
  wire xor_107473;
  wire [24:0] wide_x_squeezed;
  wire [24:0] bit_slice_107475;
  wire [27:0] shrl_107476;
  wire sticky;
  wire is_operand_inf;
  wire and_107506;
  wire is_result_nan;
  wire not_107508;
  wire p0_data_enable;
  wire bit_slice_107413;
  wire [22:0] b_fraction__6;
  wire [22:0] tuple_index_107415;
  wire [7:0] bit_slice_107416;
  wire not_107418;
  wire tuple_index_107419;
  wire [31:0] __xls_float_ips__result_buf;
  assign xls_float_ips__result_valid_inv = ~__xls_float_ips__result_valid_reg;
  assign xls_float_ips__result_valid_load_en = xls_float_ips__result_rdy | xls_float_ips__result_valid_inv;
  assign xls_float_ips__result_load_en = p7_valid & xls_float_ips__result_valid_load_en;
  assign p8_stage_done = p7_valid & xls_float_ips__result_load_en;
  assign p8_not_valid = ~p7_valid;
  assign p7_enable = p8_stage_done | p8_not_valid;
  assign p7_data_enable = p7_enable & p6_valid;
  assign p7_not_valid = ~p6_valid;
  assign p6_enable = p7_data_enable | p7_not_valid;
  assign p6_data_enable = p6_enable & p5_valid;
  assign p6_not_valid = ~p5_valid;
  assign p5_enable = p6_data_enable | p6_not_valid;
  assign p5_data_enable = p5_enable & p4_valid;
  assign p5_not_valid = ~p4_valid;
  assign p4_enable = p5_data_enable | p5_not_valid;
  assign p4_data_enable = p4_enable & p3_valid;
  assign p4_not_valid = ~p3_valid;
  assign fraction_shift__3 = 3'h4;
  assign p3_enable = p4_data_enable | p4_not_valid;
  assign add_107856 = p5_concat_107829 + 10'h001;
  assign concat_107817 = {1'h0, p4_bit_slice_107789};
  assign carry_bit = p2_abs_fraction__1[27];
  assign addend_x__2_squeezed = p1_xor_107473 ? p1_bit_slice_107475 : p1_wide_x_squeezed;
  assign a_bexp__4 = p0_bit_slice_107413 ? p0_a_bexp__2 : p0_b_bexp__6;
  assign incremented_sum__1 = p0_bit_slice_107416 + 8'h01;
  assign MAX_EXPONENT = 8'hff;
  assign a_fraction__1 = p0_bit_slice_107413 ? p0_tuple_index_107415 : p0_b_fraction__6;
  assign b_bexp__7 = p0_bit_slice_107413 ? p0_b_bexp__6 : p0_a_bexp__2;
  assign MAX_EXPONENT__1 = 8'hff;
  assign b_fraction__7 = p0_bit_slice_107413 ? p0_b_fraction__6 : p0_tuple_index_107415;
  assign p3_data_enable = p3_enable & p2_valid;
  assign p3_not_valid = ~p2_valid;
  assign wide_exponent = add_107856 - {5'h00, p5_leading_zeroes__4_to_5, p5_leading_zeroes__0_to_4};
  assign do_round_up = p4_normal_chunk > fraction_shift__3 | p4_half_way_chunk == 2'h3;
  assign add_107820 = concat_107817 + 25'h000_0001;
  assign leading_zeroes__0_to_4 = priority_sel_4b_2way({p3_nor_107730, p3_leading_zeroes__4_to_5}, {p3_and_107697, p3_priority_sel_107732}, {1'h1, p3_nor_107703, p3_priority_sel_107733}, {p3_and_107695, p3_priority_sel_107734});
  assign nor_107602 = ~(p2_abs_fraction__1[11] | p2_abs_fraction__1[10]);
  assign nor_107603 = ~(p2_abs_fraction__1[9] | p2_abs_fraction__1[8]);
  assign nor_107605 = ~(p2_abs_fraction__1[1] | p2_abs_fraction__1[0]);
  assign nor_107606 = ~(p2_abs_fraction__1[3] | p2_abs_fraction__1[2]);
  assign nor_107611 = ~(p2_abs_fraction__1[5] | p2_abs_fraction__1[4]);
  assign nor_107612 = ~(p2_abs_fraction__1[7] | p2_abs_fraction__1[6]);
  assign nor_107617 = ~(p2_abs_fraction__1[17] | p2_abs_fraction__1[16]);
  assign nor_107620 = ~(p2_abs_fraction__1[13] | p2_abs_fraction__1[12]);
  assign nor_107621 = ~(carry_bit | p2_abs_fraction__1[26]);
  assign nor_107622 = ~(p2_abs_fraction__1[25] | p2_abs_fraction__1[24]);
  assign nor_107628 = ~(p2_abs_fraction__1[21] | p2_abs_fraction__1[20]);
  assign a_bexpbs_difference__2 = p0_bit_slice_107413 ? incremented_sum__1 : ~p0_bit_slice_107416;
  assign eq_107486 = a_bexp__4 == MAX_EXPONENT;
  assign eq_107487 = a_fraction__1 == 23'h00_0000;
  assign eq_107488 = b_bexp__7 == MAX_EXPONENT__1;
  assign eq_107489 = b_fraction__7 == 23'h00_0000;
  assign p2_enable = p3_data_enable | p3_not_valid;
  assign and_reduce_107883 = &p6_wide_exponent__2[7:0];
  assign wide_exponent__1 = wide_exponent & {10{p5_not_107554}};
  assign rounded_fraction_squeezed_portion_3_width_25 = do_round_up ? add_107820 : concat_107817;
  assign leading_zeroes = {p3_leading_zeroes__4_to_5, leading_zeroes__0_to_4};
  assign nor_107629 = ~(p2_abs_fraction__1[23] | p2_abs_fraction__1[22]);
  assign and_107630 = nor_107602 & nor_107603;
  assign and_107632 = nor_107606 & nor_107605;
  assign nor_107637 = ~(p2_abs_fraction__1[7] | p2_abs_fraction__1[6] | nor_107611);
  assign and_107638 = nor_107612 & nor_107611;
  assign nor_107641 = ~(p2_abs_fraction__1[11] | ~p2_abs_fraction__1[10]);
  assign and_107645 = ~(p2_abs_fraction__1[19] | p2_abs_fraction__1[18]) & nor_107617;
  assign nor_107646 = ~(p2_abs_fraction__1[15] | p2_abs_fraction__1[14]);
  assign and_107650 = nor_107621 & nor_107622;
  assign nor_107652 = ~(carry_bit | ~p2_abs_fraction__1[26]);
  assign add_107538 = {{1{addend_x__2_squeezed[24]}}, addend_x__2_squeezed} + {1'h0, p1_shrl_107476[27:3]};
  assign fraction_x = {1'h1, a_fraction__1};
  assign a_sign__1 = p0_bit_slice_107413 ? p0_tuple_index_107419 : p0_not_107418;
  assign b_sign__3 = p0_bit_slice_107413 ? p0_not_107418 : p0_tuple_index_107419;
  assign p2_data_enable = p2_enable & p1_valid;
  assign p2_not_valid = ~p1_valid;
  assign b_bexp__6 = xls_float_ips__rhs[30:23];
  assign rounding_carry = rounded_fraction_squeezed_portion_3_width_25[24];
  assign fraction_shift__2 = 3'h3;
  assign fraction_shift__4 = 3'h4;
  assign cancel_fraction = leading_zeroes >= 5'h1d ? 29'h0000_0000 : {1'h0, p3_abs_fraction__1} << leading_zeroes;
  assign and_107659 = nor_107629 & nor_107628;
  assign and_107677 = nor_107646 & nor_107620;
  assign fraction_x__1 = fraction_x & {24{a_bexp__4 != 8'h00}};
  assign addend_x__2_squeezed_const_lsb_bits__1 = 3'h0;
  assign fraction_y = {1'h1, b_fraction__7};
  assign sign_ext_107458 = {24{b_bexp__7 != 8'h00}};
  assign add_107477 = (a_bexpbs_difference__2 >= 8'h1c ? 28'h000_0000 : 28'h000_0001 << a_bexpbs_difference__2) + 28'hfff_ffff;
  assign p1_enable = p2_data_enable | p2_not_valid;
  assign a_bexp__2 = xls_float_ips__lhs[30:23];
  assign rounded_fraction = {rounded_fraction_squeezed_portion_3_width_25, p4_normal_chunk};
  assign fraction_shift__1 = rounding_carry ? fraction_shift__4 : fraction_shift__2;
  assign cancel_fraction__1 = cancel_fraction[27:1];
  assign carry_fraction__1 = {p3_abs_fraction__1[27:2], p3_or_107735};
  assign and_107695 = and_107650 & and_107659;
  assign and_107697 = and_107630 & and_107638;
  assign nor_107703 = ~(~and_107645 | and_107677);
  assign and_107704 = and_107645 & and_107677;
  assign priority_sel_107711 = priority_sel_2b_2way({~(carry_bit | p2_abs_fraction__1[26] | nor_107622), and_107650}, {nor_107652, 1'h0}, {1'h1, ~(p2_abs_fraction__1[25] | ~p2_abs_fraction__1[24])}, {nor_107621, nor_107652});
  assign concat_107543 = {add_107538[24:0], p1_shrl_107476[2:1], p1_shrl_107476[0] | p1_sticky};
  assign fraction_is_zero = add_107538 == 26'h000_0000 & ~(p1_shrl_107476[1] | p1_shrl_107476[2]) & ~(p1_shrl_107476[0] | p1_sticky);
  assign wide_x = {1'h0, fraction_x__1, addend_x__2_squeezed_const_lsb_bits__1};
  assign fraction_y__1 = fraction_y & sign_ext_107458;
  assign addend_x__2_squeezed_const_lsb_bits = 3'h0;
  assign has_pos_inf = ~(~eq_107486 | ~eq_107487 | a_sign__1) | ~(~eq_107488 | ~eq_107489 | b_sign__3);
  assign has_neg_inf = eq_107486 & eq_107487 & a_sign__1 | eq_107488 & eq_107489 & b_sign__3;
  assign p1_data_enable = p1_enable & p0_valid;
  assign p1_not_valid = ~p0_valid;
  assign FRACTION_HIGH_BIT = 23'h40_0000;
  assign sign_ext_107887 = {23{~(p6_is_operand_inf | p6_wide_exponent__2[8] | and_reduce_107883 | ~((|p6_wide_exponent__2[8:1]) | p6_wide_exponent__2[0]))}};
  assign MAX_EXPONENT__2 = 8'hff;
  assign add_107828 = {1'h0, p4_a_bexp__4} + {8'h00, rounding_carry};
  assign shrl_107834 = rounded_fraction >> fraction_shift__1;
  assign shifted_fraction = p3_carry_bit ? carry_fraction__1 : cancel_fraction__1;
  assign concat_107717 = {and_107632, priority_sel_2b_2way({~(p2_abs_fraction__1[3] | p2_abs_fraction__1[2] | nor_107605), and_107632}, 2'h0, {1'h1, ~(p2_abs_fraction__1[1] | ~p2_abs_fraction__1[0])}, {nor_107606, ~(p2_abs_fraction__1[3] | ~p2_abs_fraction__1[2])})};
  assign concat_107718 = {1'h1, nor_107637, priority_sel_1b_4way({~(p2_abs_fraction__1[7] | ~p2_abs_fraction__1[6]), nor_107612, nor_107637, and_107638}, 1'h0, ~(p2_abs_fraction__1[5] | ~p2_abs_fraction__1[4]), 1'h0, 1'h1, 1'h0)};
  assign concat_107719 = {and_107630, priority_sel_2b_2way({~(p2_abs_fraction__1[11] | p2_abs_fraction__1[10] | nor_107603), and_107630}, {nor_107641, 1'h0}, {1'h1, ~(p2_abs_fraction__1[9] | ~p2_abs_fraction__1[8])}, {nor_107602, nor_107641})};
  assign concat_107722 = {nor_107646, priority_sel_1b_3way({~(p2_abs_fraction__1[15] | ~p2_abs_fraction__1[14]), nor_107646, ~(p2_abs_fraction__1[15] | p2_abs_fraction__1[14] | nor_107620)}, ~(p2_abs_fraction__1[13] | ~p2_abs_fraction__1[12]), 1'h0, 1'h1, 1'h0)};
  assign concat_107728 = {1'h1, nor_107629, priority_sel_1b_3way({~(p2_abs_fraction__1[23] | ~p2_abs_fraction__1[22]), nor_107629, ~(p2_abs_fraction__1[23] | p2_abs_fraction__1[22] | nor_107628)}, ~(p2_abs_fraction__1[21] | ~p2_abs_fraction__1[20]), 1'h0, 1'h1, 1'h0)};
  assign result_sign__1 = p2_is_operand_inf ? p2_not_107508 : p2_result_sign;
  assign neg_107469 = -wide_x;
  assign wide_y = {1'h0, fraction_y__1, addend_x__2_squeezed_const_lsb_bits};
  assign p0_enable = p1_data_enable | p1_not_valid;
  assign p0_all_active_inputs_valid = xls_float_ips__rhs_vld & xls_float_ips__lhs_vld;
  assign sum = {1'h0, a_bexp__2} + {1'h0, ~b_bexp__6};
  assign b_sign__2 = xls_float_ips__rhs[31:31];
  assign result_fraction__4 = p7_is_result_nan ? FRACTION_HIGH_BIT : p7_result_fraction__3;
  assign result_fraction__3 = p6_result_fraction & sign_ext_107887;
  assign result_exponent__2 = p6_is_result_nan | p6_is_operand_inf | p6_wide_exponent__2[8] | and_reduce_107883 ? MAX_EXPONENT__2 : p6_wide_exponent__2[7:0];
  assign wide_exponent__2 = wide_exponent__1[8:0] & {9{~wide_exponent__1[9]}};
  assign concat_107829 = {1'h0, add_107828};
  assign result_fraction = shrl_107834[22:0];
  assign normal_chunk = shifted_fraction[2:0];
  assign half_way_chunk = shifted_fraction[3:2];
  assign bit_slice_107789 = shifted_fraction[26:3];
  assign nor_107730 = ~(~and_107695 | and_107704);
  assign leading_zeroes__4_to_5 = and_107695 & and_107704;
  assign priority_sel_107732 = priority_sel_3b_2way({~(~and_107630 | and_107638), and_107697}, concat_107717, concat_107718, concat_107719);
  assign priority_sel_107733 = priority_sel_2b_4way({~(p2_abs_fraction__1[19] | p2_abs_fraction__1[18] | nor_107617), and_107645, nor_107703, and_107704}, 2'h0, concat_107722, 2'h0, {1'h1, ~(p2_abs_fraction__1[17] | ~p2_abs_fraction__1[16])}, {1'h0, ~(p2_abs_fraction__1[19] | ~p2_abs_fraction__1[18])});
  assign priority_sel_107734 = priority_sel_3b_2way({~(~and_107650 | and_107659), and_107695}, {priority_sel_107711, 1'h0}, concat_107728, {and_107650, priority_sel_107711});
  assign or_107735 = p2_abs_fraction__1[1] | p2_abs_fraction__1[0];
  assign result_sign__2 = ~p2_is_result_nan & result_sign__1;
  assign abs_fraction__1 = add_107538[25] ? -concat_107543 : concat_107543;
  assign not_107554 = ~fraction_is_zero;
  assign result_sign = priority_sel_1b_2way({add_107538[25], fraction_is_zero}, p1_and_107506, ~p1_b_sign__3, p1_b_sign__3);
  assign xor_107473 = a_sign__1 ^ b_sign__3;
  assign wide_x_squeezed = {1'h0, fraction_x__1};
  assign bit_slice_107475 = neg_107469[27:3];
  assign shrl_107476 = a_bexpbs_difference__2 >= 8'h1c ? 28'h000_0000 : wide_y >> a_bexpbs_difference__2;
  assign sticky = (fraction_y & sign_ext_107458 & add_107477[26:3]) != 24'h00_0000;
  assign is_operand_inf = eq_107486 & eq_107487 | eq_107488 & eq_107489;
  assign and_107506 = a_sign__1 & b_sign__3;
  assign is_result_nan = ~(~eq_107486 | eq_107487) | ~(~eq_107488 | eq_107489) | has_pos_inf & has_neg_inf;
  assign not_107508 = ~has_pos_inf;
  assign p0_data_enable = p0_enable & p0_all_active_inputs_valid;
  assign bit_slice_107413 = sum[8];
  assign b_fraction__6 = xls_float_ips__rhs[22:0];
  assign tuple_index_107415 = xls_float_ips__lhs[22:0];
  assign bit_slice_107416 = sum[7:0];
  assign not_107418 = ~b_sign__2;
  assign tuple_index_107419 = xls_float_ips__lhs[31:31];
  assign __xls_float_ips__result_buf = {p7_result_sign__2, p7_result_exponent__2, result_fraction__4};
  always @ (posedge clk) begin
    if (rst) begin
      p0_b_bexp__6 <= 8'h00;
      p0_a_bexp__2 <= 8'h00;
      p0_bit_slice_107413 <= 1'h0;
      p0_b_fraction__6 <= 23'h00_0000;
      p0_tuple_index_107415 <= 23'h00_0000;
      p0_bit_slice_107416 <= 8'h00;
      p0_not_107418 <= 1'h0;
      p0_tuple_index_107419 <= 1'h0;
      p1_a_bexp__4 <= 8'h00;
      p1_b_sign__3 <= 1'h0;
      p1_xor_107473 <= 1'h0;
      p1_wide_x_squeezed <= 25'h000_0000;
      p1_bit_slice_107475 <= 25'h000_0000;
      p1_shrl_107476 <= 28'h000_0000;
      p1_sticky <= 1'h0;
      p1_is_operand_inf <= 1'h0;
      p1_and_107506 <= 1'h0;
      p1_is_result_nan <= 1'h0;
      p1_not_107508 <= 1'h0;
      p2_a_bexp__4 <= 8'h00;
      p2_abs_fraction__1 <= 28'h000_0000;
      p2_not_107554 <= 1'h0;
      p2_is_operand_inf <= 1'h0;
      p2_is_result_nan <= 1'h0;
      p2_result_sign <= 1'h0;
      p2_not_107508 <= 1'h0;
      p3_a_bexp__4 <= 8'h00;
      p3_abs_fraction__1 <= 28'h000_0000;
      p3_carry_bit <= 1'h0;
      p3_and_107695 <= 1'h0;
      p3_and_107697 <= 1'h0;
      p3_nor_107703 <= 1'h0;
      p3_nor_107730 <= 1'h0;
      p3_leading_zeroes__4_to_5 <= 1'h0;
      p3_priority_sel_107732 <= 3'h0;
      p3_priority_sel_107733 <= 2'h0;
      p3_priority_sel_107734 <= 3'h0;
      p3_or_107735 <= 1'h0;
      p3_not_107554 <= 1'h0;
      p3_is_operand_inf <= 1'h0;
      p3_is_result_nan <= 1'h0;
      p3_result_sign__2 <= 1'h0;
      p4_a_bexp__4 <= 8'h00;
      p4_leading_zeroes__4_to_5 <= 1'h0;
      p4_leading_zeroes__0_to_4 <= 4'h0;
      p4_normal_chunk <= 3'h0;
      p4_half_way_chunk <= 2'h0;
      p4_bit_slice_107789 <= 24'h00_0000;
      p4_not_107554 <= 1'h0;
      p4_is_operand_inf <= 1'h0;
      p4_is_result_nan <= 1'h0;
      p4_result_sign__2 <= 1'h0;
      p5_leading_zeroes__4_to_5 <= 1'h0;
      p5_leading_zeroes__0_to_4 <= 4'h0;
      p5_concat_107829 <= 10'h000;
      p5_not_107554 <= 1'h0;
      p5_is_operand_inf <= 1'h0;
      p5_is_result_nan <= 1'h0;
      p5_result_fraction <= 23'h00_0000;
      p5_result_sign__2 <= 1'h0;
      p6_wide_exponent__2 <= 9'h000;
      p6_is_operand_inf <= 1'h0;
      p6_is_result_nan <= 1'h0;
      p6_result_fraction <= 23'h00_0000;
      p6_result_sign__2 <= 1'h0;
      p7_is_result_nan <= 1'h0;
      p7_result_fraction__3 <= 23'h00_0000;
      p7_result_sign__2 <= 1'h0;
      p7_result_exponent__2 <= 8'h00;
      p0_valid <= 1'h0;
      p1_valid <= 1'h0;
      p2_valid <= 1'h0;
      p3_valid <= 1'h0;
      p4_valid <= 1'h0;
      p5_valid <= 1'h0;
      p6_valid <= 1'h0;
      p7_valid <= 1'h0;
      __xls_float_ips__result_reg <= __xls_float_ips__result_reg_init;
      __xls_float_ips__result_valid_reg <= 1'h0;
    end else begin
      p0_b_bexp__6 <= p0_data_enable ? b_bexp__6 : p0_b_bexp__6;
      p0_a_bexp__2 <= p0_data_enable ? a_bexp__2 : p0_a_bexp__2;
      p0_bit_slice_107413 <= p0_data_enable ? bit_slice_107413 : p0_bit_slice_107413;
      p0_b_fraction__6 <= p0_data_enable ? b_fraction__6 : p0_b_fraction__6;
      p0_tuple_index_107415 <= p0_data_enable ? tuple_index_107415 : p0_tuple_index_107415;
      p0_bit_slice_107416 <= p0_data_enable ? bit_slice_107416 : p0_bit_slice_107416;
      p0_not_107418 <= p0_data_enable ? not_107418 : p0_not_107418;
      p0_tuple_index_107419 <= p0_data_enable ? tuple_index_107419 : p0_tuple_index_107419;
      p1_a_bexp__4 <= p1_data_enable ? a_bexp__4 : p1_a_bexp__4;
      p1_b_sign__3 <= p1_data_enable ? b_sign__3 : p1_b_sign__3;
      p1_xor_107473 <= p1_data_enable ? xor_107473 : p1_xor_107473;
      p1_wide_x_squeezed <= p1_data_enable ? wide_x_squeezed : p1_wide_x_squeezed;
      p1_bit_slice_107475 <= p1_data_enable ? bit_slice_107475 : p1_bit_slice_107475;
      p1_shrl_107476 <= p1_data_enable ? shrl_107476 : p1_shrl_107476;
      p1_sticky <= p1_data_enable ? sticky : p1_sticky;
      p1_is_operand_inf <= p1_data_enable ? is_operand_inf : p1_is_operand_inf;
      p1_and_107506 <= p1_data_enable ? and_107506 : p1_and_107506;
      p1_is_result_nan <= p1_data_enable ? is_result_nan : p1_is_result_nan;
      p1_not_107508 <= p1_data_enable ? not_107508 : p1_not_107508;
      p2_a_bexp__4 <= p2_data_enable ? p1_a_bexp__4 : p2_a_bexp__4;
      p2_abs_fraction__1 <= p2_data_enable ? abs_fraction__1 : p2_abs_fraction__1;
      p2_not_107554 <= p2_data_enable ? not_107554 : p2_not_107554;
      p2_is_operand_inf <= p2_data_enable ? p1_is_operand_inf : p2_is_operand_inf;
      p2_is_result_nan <= p2_data_enable ? p1_is_result_nan : p2_is_result_nan;
      p2_result_sign <= p2_data_enable ? result_sign : p2_result_sign;
      p2_not_107508 <= p2_data_enable ? p1_not_107508 : p2_not_107508;
      p3_a_bexp__4 <= p3_data_enable ? p2_a_bexp__4 : p3_a_bexp__4;
      p3_abs_fraction__1 <= p3_data_enable ? p2_abs_fraction__1 : p3_abs_fraction__1;
      p3_carry_bit <= p3_data_enable ? carry_bit : p3_carry_bit;
      p3_and_107695 <= p3_data_enable ? and_107695 : p3_and_107695;
      p3_and_107697 <= p3_data_enable ? and_107697 : p3_and_107697;
      p3_nor_107703 <= p3_data_enable ? nor_107703 : p3_nor_107703;
      p3_nor_107730 <= p3_data_enable ? nor_107730 : p3_nor_107730;
      p3_leading_zeroes__4_to_5 <= p3_data_enable ? leading_zeroes__4_to_5 : p3_leading_zeroes__4_to_5;
      p3_priority_sel_107732 <= p3_data_enable ? priority_sel_107732 : p3_priority_sel_107732;
      p3_priority_sel_107733 <= p3_data_enable ? priority_sel_107733 : p3_priority_sel_107733;
      p3_priority_sel_107734 <= p3_data_enable ? priority_sel_107734 : p3_priority_sel_107734;
      p3_or_107735 <= p3_data_enable ? or_107735 : p3_or_107735;
      p3_not_107554 <= p3_data_enable ? p2_not_107554 : p3_not_107554;
      p3_is_operand_inf <= p3_data_enable ? p2_is_operand_inf : p3_is_operand_inf;
      p3_is_result_nan <= p3_data_enable ? p2_is_result_nan : p3_is_result_nan;
      p3_result_sign__2 <= p3_data_enable ? result_sign__2 : p3_result_sign__2;
      p4_a_bexp__4 <= p4_data_enable ? p3_a_bexp__4 : p4_a_bexp__4;
      p4_leading_zeroes__4_to_5 <= p4_data_enable ? p3_leading_zeroes__4_to_5 : p4_leading_zeroes__4_to_5;
      p4_leading_zeroes__0_to_4 <= p4_data_enable ? leading_zeroes__0_to_4 : p4_leading_zeroes__0_to_4;
      p4_normal_chunk <= p4_data_enable ? normal_chunk : p4_normal_chunk;
      p4_half_way_chunk <= p4_data_enable ? half_way_chunk : p4_half_way_chunk;
      p4_bit_slice_107789 <= p4_data_enable ? bit_slice_107789 : p4_bit_slice_107789;
      p4_not_107554 <= p4_data_enable ? p3_not_107554 : p4_not_107554;
      p4_is_operand_inf <= p4_data_enable ? p3_is_operand_inf : p4_is_operand_inf;
      p4_is_result_nan <= p4_data_enable ? p3_is_result_nan : p4_is_result_nan;
      p4_result_sign__2 <= p4_data_enable ? p3_result_sign__2 : p4_result_sign__2;
      p5_leading_zeroes__4_to_5 <= p5_data_enable ? p4_leading_zeroes__4_to_5 : p5_leading_zeroes__4_to_5;
      p5_leading_zeroes__0_to_4 <= p5_data_enable ? p4_leading_zeroes__0_to_4 : p5_leading_zeroes__0_to_4;
      p5_concat_107829 <= p5_data_enable ? concat_107829 : p5_concat_107829;
      p5_not_107554 <= p5_data_enable ? p4_not_107554 : p5_not_107554;
      p5_is_operand_inf <= p5_data_enable ? p4_is_operand_inf : p5_is_operand_inf;
      p5_is_result_nan <= p5_data_enable ? p4_is_result_nan : p5_is_result_nan;
      p5_result_fraction <= p5_data_enable ? result_fraction : p5_result_fraction;
      p5_result_sign__2 <= p5_data_enable ? p4_result_sign__2 : p5_result_sign__2;
      p6_wide_exponent__2 <= p6_data_enable ? wide_exponent__2 : p6_wide_exponent__2;
      p6_is_operand_inf <= p6_data_enable ? p5_is_operand_inf : p6_is_operand_inf;
      p6_is_result_nan <= p6_data_enable ? p5_is_result_nan : p6_is_result_nan;
      p6_result_fraction <= p6_data_enable ? p5_result_fraction : p6_result_fraction;
      p6_result_sign__2 <= p6_data_enable ? p5_result_sign__2 : p6_result_sign__2;
      p7_is_result_nan <= p7_data_enable ? p6_is_result_nan : p7_is_result_nan;
      p7_result_fraction__3 <= p7_data_enable ? result_fraction__3 : p7_result_fraction__3;
      p7_result_sign__2 <= p7_data_enable ? p6_result_sign__2 : p7_result_sign__2;
      p7_result_exponent__2 <= p7_data_enable ? result_exponent__2 : p7_result_exponent__2;
      p0_valid <= p0_enable ? p0_all_active_inputs_valid : p0_valid;
      p1_valid <= p1_enable ? p0_valid : p1_valid;
      p2_valid <= p2_enable ? p1_valid : p2_valid;
      p3_valid <= p3_enable ? p2_valid : p3_valid;
      p4_valid <= p4_enable ? p3_valid : p4_valid;
      p5_valid <= p5_enable ? p4_valid : p5_valid;
      p6_valid <= p6_enable ? p5_valid : p6_valid;
      p7_valid <= p7_enable ? p6_valid : p7_valid;
      __xls_float_ips__result_reg <= xls_float_ips__result_load_en ? __xls_float_ips__result_buf : __xls_float_ips__result_reg;
      __xls_float_ips__result_valid_reg <= xls_float_ips__result_valid_load_en ? p7_valid : __xls_float_ips__result_valid_reg;
    end
  end
  assign xls_float_ips__result = __xls_float_ips__result_reg;
  assign xls_float_ips__result_vld = __xls_float_ips__result_valid_reg;
  assign xls_float_ips__rhs_rdy = p0_data_enable;
  assign xls_float_ips__lhs_rdy = p0_data_enable;
endmodule
