library ieee;
use ieee.std_logic_1164.all;

package types is
  type data_array is array(natural range <>) of std_logic_vector;
end package;
